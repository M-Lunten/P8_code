-- megafunction wizard: %LPM_MUX%
-- GENERATION: STANDARD
-- VERSION: WM1.0
-- MODULE: LPM_MUX 

-- ============================================================
-- File Name: out_mux.vhd
-- Megafunction Name(s):
-- 			LPM_MUX
--
-- Simulation Library Files(s):
-- 			lpm
-- ============================================================
-- ************************************************************
-- THIS IS A WIZARD-GENERATED FILE. DO NOT EDIT THIS FILE!
--
-- 18.1.0 Build 625 09/12/2018 SJ Lite Edition
-- ************************************************************


--Copyright (C) 2018  Intel Corporation. All rights reserved.
--Your use of Intel Corporation's design tools, logic functions 
--and other software and tools, and its AMPP partner logic 
--functions, and any output files from any of the foregoing 
--(including device programming or simulation files), and any 
--associated documentation or information are expressly subject 
--to the terms and conditions of the Intel Program License 
--Subscription Agreement, the Intel Quartus Prime License Agreement,
--the Intel FPGA IP License Agreement, or other applicable license
--agreement, including, without limitation, that your use is for
--the sole purpose of programming logic devices manufactured by
--Intel and sold by Intel or its authorized distributors.  Please
--refer to the applicable agreement for further details.


LIBRARY ieee;
USE ieee.std_logic_1164.all;

LIBRARY lpm;
USE lpm.lpm_components.all;

ENTITY out_mux IS
	PORT
	(
		data0x		: IN STD_LOGIC_VECTOR (31 DOWNTO 0);
		data100x		: IN STD_LOGIC_VECTOR (31 DOWNTO 0);
		data101x		: IN STD_LOGIC_VECTOR (31 DOWNTO 0);
		data102x		: IN STD_LOGIC_VECTOR (31 DOWNTO 0);
		data103x		: IN STD_LOGIC_VECTOR (31 DOWNTO 0);
		data104x		: IN STD_LOGIC_VECTOR (31 DOWNTO 0);
		data105x		: IN STD_LOGIC_VECTOR (31 DOWNTO 0);
		data106x		: IN STD_LOGIC_VECTOR (31 DOWNTO 0);
		data107x		: IN STD_LOGIC_VECTOR (31 DOWNTO 0);
		data108x		: IN STD_LOGIC_VECTOR (31 DOWNTO 0);
		data109x		: IN STD_LOGIC_VECTOR (31 DOWNTO 0);
		data10x		: IN STD_LOGIC_VECTOR (31 DOWNTO 0);
		data110x		: IN STD_LOGIC_VECTOR (31 DOWNTO 0);
		data111x		: IN STD_LOGIC_VECTOR (31 DOWNTO 0);
		data112x		: IN STD_LOGIC_VECTOR (31 DOWNTO 0);
		data113x		: IN STD_LOGIC_VECTOR (31 DOWNTO 0);
		data114x		: IN STD_LOGIC_VECTOR (31 DOWNTO 0);
		data115x		: IN STD_LOGIC_VECTOR (31 DOWNTO 0);
		data116x		: IN STD_LOGIC_VECTOR (31 DOWNTO 0);
		data117x		: IN STD_LOGIC_VECTOR (31 DOWNTO 0);
		data118x		: IN STD_LOGIC_VECTOR (31 DOWNTO 0);
		data119x		: IN STD_LOGIC_VECTOR (31 DOWNTO 0);
		data11x		: IN STD_LOGIC_VECTOR (31 DOWNTO 0);
		data120x		: IN STD_LOGIC_VECTOR (31 DOWNTO 0);
		data121x		: IN STD_LOGIC_VECTOR (31 DOWNTO 0);
		data122x		: IN STD_LOGIC_VECTOR (31 DOWNTO 0);
		data123x		: IN STD_LOGIC_VECTOR (31 DOWNTO 0);
		data124x		: IN STD_LOGIC_VECTOR (31 DOWNTO 0);
		data125x		: IN STD_LOGIC_VECTOR (31 DOWNTO 0);
		data126x		: IN STD_LOGIC_VECTOR (31 DOWNTO 0);
		data127x		: IN STD_LOGIC_VECTOR (31 DOWNTO 0);
		data12x		: IN STD_LOGIC_VECTOR (31 DOWNTO 0);
		data13x		: IN STD_LOGIC_VECTOR (31 DOWNTO 0);
		data14x		: IN STD_LOGIC_VECTOR (31 DOWNTO 0);
		data15x		: IN STD_LOGIC_VECTOR (31 DOWNTO 0);
		data16x		: IN STD_LOGIC_VECTOR (31 DOWNTO 0);
		data17x		: IN STD_LOGIC_VECTOR (31 DOWNTO 0);
		data18x		: IN STD_LOGIC_VECTOR (31 DOWNTO 0);
		data19x		: IN STD_LOGIC_VECTOR (31 DOWNTO 0);
		data1x		: IN STD_LOGIC_VECTOR (31 DOWNTO 0);
		data20x		: IN STD_LOGIC_VECTOR (31 DOWNTO 0);
		data21x		: IN STD_LOGIC_VECTOR (31 DOWNTO 0);
		data22x		: IN STD_LOGIC_VECTOR (31 DOWNTO 0);
		data23x		: IN STD_LOGIC_VECTOR (31 DOWNTO 0);
		data24x		: IN STD_LOGIC_VECTOR (31 DOWNTO 0);
		data25x		: IN STD_LOGIC_VECTOR (31 DOWNTO 0);
		data26x		: IN STD_LOGIC_VECTOR (31 DOWNTO 0);
		data27x		: IN STD_LOGIC_VECTOR (31 DOWNTO 0);
		data28x		: IN STD_LOGIC_VECTOR (31 DOWNTO 0);
		data29x		: IN STD_LOGIC_VECTOR (31 DOWNTO 0);
		data2x		: IN STD_LOGIC_VECTOR (31 DOWNTO 0);
		data30x		: IN STD_LOGIC_VECTOR (31 DOWNTO 0);
		data31x		: IN STD_LOGIC_VECTOR (31 DOWNTO 0);
		data32x		: IN STD_LOGIC_VECTOR (31 DOWNTO 0);
		data33x		: IN STD_LOGIC_VECTOR (31 DOWNTO 0);
		data34x		: IN STD_LOGIC_VECTOR (31 DOWNTO 0);
		data35x		: IN STD_LOGIC_VECTOR (31 DOWNTO 0);
		data36x		: IN STD_LOGIC_VECTOR (31 DOWNTO 0);
		data37x		: IN STD_LOGIC_VECTOR (31 DOWNTO 0);
		data38x		: IN STD_LOGIC_VECTOR (31 DOWNTO 0);
		data39x		: IN STD_LOGIC_VECTOR (31 DOWNTO 0);
		data3x		: IN STD_LOGIC_VECTOR (31 DOWNTO 0);
		data40x		: IN STD_LOGIC_VECTOR (31 DOWNTO 0);
		data41x		: IN STD_LOGIC_VECTOR (31 DOWNTO 0);
		data42x		: IN STD_LOGIC_VECTOR (31 DOWNTO 0);
		data43x		: IN STD_LOGIC_VECTOR (31 DOWNTO 0);
		data44x		: IN STD_LOGIC_VECTOR (31 DOWNTO 0);
		data45x		: IN STD_LOGIC_VECTOR (31 DOWNTO 0);
		data46x		: IN STD_LOGIC_VECTOR (31 DOWNTO 0);
		data47x		: IN STD_LOGIC_VECTOR (31 DOWNTO 0);
		data48x		: IN STD_LOGIC_VECTOR (31 DOWNTO 0);
		data49x		: IN STD_LOGIC_VECTOR (31 DOWNTO 0);
		data4x		: IN STD_LOGIC_VECTOR (31 DOWNTO 0);
		data50x		: IN STD_LOGIC_VECTOR (31 DOWNTO 0);
		data51x		: IN STD_LOGIC_VECTOR (31 DOWNTO 0);
		data52x		: IN STD_LOGIC_VECTOR (31 DOWNTO 0);
		data53x		: IN STD_LOGIC_VECTOR (31 DOWNTO 0);
		data54x		: IN STD_LOGIC_VECTOR (31 DOWNTO 0);
		data55x		: IN STD_LOGIC_VECTOR (31 DOWNTO 0);
		data56x		: IN STD_LOGIC_VECTOR (31 DOWNTO 0);
		data57x		: IN STD_LOGIC_VECTOR (31 DOWNTO 0);
		data58x		: IN STD_LOGIC_VECTOR (31 DOWNTO 0);
		data59x		: IN STD_LOGIC_VECTOR (31 DOWNTO 0);
		data5x		: IN STD_LOGIC_VECTOR (31 DOWNTO 0);
		data60x		: IN STD_LOGIC_VECTOR (31 DOWNTO 0);
		data61x		: IN STD_LOGIC_VECTOR (31 DOWNTO 0);
		data62x		: IN STD_LOGIC_VECTOR (31 DOWNTO 0);
		data63x		: IN STD_LOGIC_VECTOR (31 DOWNTO 0);
		data64x		: IN STD_LOGIC_VECTOR (31 DOWNTO 0);
		data65x		: IN STD_LOGIC_VECTOR (31 DOWNTO 0);
		data66x		: IN STD_LOGIC_VECTOR (31 DOWNTO 0);
		data67x		: IN STD_LOGIC_VECTOR (31 DOWNTO 0);
		data68x		: IN STD_LOGIC_VECTOR (31 DOWNTO 0);
		data69x		: IN STD_LOGIC_VECTOR (31 DOWNTO 0);
		data6x		: IN STD_LOGIC_VECTOR (31 DOWNTO 0);
		data70x		: IN STD_LOGIC_VECTOR (31 DOWNTO 0);
		data71x		: IN STD_LOGIC_VECTOR (31 DOWNTO 0);
		data72x		: IN STD_LOGIC_VECTOR (31 DOWNTO 0);
		data73x		: IN STD_LOGIC_VECTOR (31 DOWNTO 0);
		data74x		: IN STD_LOGIC_VECTOR (31 DOWNTO 0);
		data75x		: IN STD_LOGIC_VECTOR (31 DOWNTO 0);
		data76x		: IN STD_LOGIC_VECTOR (31 DOWNTO 0);
		data77x		: IN STD_LOGIC_VECTOR (31 DOWNTO 0);
		data78x		: IN STD_LOGIC_VECTOR (31 DOWNTO 0);
		data79x		: IN STD_LOGIC_VECTOR (31 DOWNTO 0);
		data7x		: IN STD_LOGIC_VECTOR (31 DOWNTO 0);
		data80x		: IN STD_LOGIC_VECTOR (31 DOWNTO 0);
		data81x		: IN STD_LOGIC_VECTOR (31 DOWNTO 0);
		data82x		: IN STD_LOGIC_VECTOR (31 DOWNTO 0);
		data83x		: IN STD_LOGIC_VECTOR (31 DOWNTO 0);
		data84x		: IN STD_LOGIC_VECTOR (31 DOWNTO 0);
		data85x		: IN STD_LOGIC_VECTOR (31 DOWNTO 0);
		data86x		: IN STD_LOGIC_VECTOR (31 DOWNTO 0);
		data87x		: IN STD_LOGIC_VECTOR (31 DOWNTO 0);
		data88x		: IN STD_LOGIC_VECTOR (31 DOWNTO 0);
		data89x		: IN STD_LOGIC_VECTOR (31 DOWNTO 0);
		data8x		: IN STD_LOGIC_VECTOR (31 DOWNTO 0);
		data90x		: IN STD_LOGIC_VECTOR (31 DOWNTO 0);
		data91x		: IN STD_LOGIC_VECTOR (31 DOWNTO 0);
		data92x		: IN STD_LOGIC_VECTOR (31 DOWNTO 0);
		data93x		: IN STD_LOGIC_VECTOR (31 DOWNTO 0);
		data94x		: IN STD_LOGIC_VECTOR (31 DOWNTO 0);
		data95x		: IN STD_LOGIC_VECTOR (31 DOWNTO 0);
		data96x		: IN STD_LOGIC_VECTOR (31 DOWNTO 0);
		data97x		: IN STD_LOGIC_VECTOR (31 DOWNTO 0);
		data98x		: IN STD_LOGIC_VECTOR (31 DOWNTO 0);
		data99x		: IN STD_LOGIC_VECTOR (31 DOWNTO 0);
		data9x		: IN STD_LOGIC_VECTOR (31 DOWNTO 0);
		sel		: IN STD_LOGIC_VECTOR (6 DOWNTO 0);
		result		: OUT STD_LOGIC_VECTOR (31 DOWNTO 0)
	);
END out_mux;


ARCHITECTURE SYN OF out_mux IS

--	type STD_LOGIC_2D is array (NATURAL RANGE <>, NATURAL RANGE <>) of STD_LOGIC;

	SIGNAL sub_wire0	: STD_LOGIC_VECTOR (31 DOWNTO 0);
	SIGNAL sub_wire1	: STD_LOGIC_2D (127 DOWNTO 0, 31 DOWNTO 0);
	SIGNAL sub_wire2	: STD_LOGIC_VECTOR (31 DOWNTO 0);
	SIGNAL sub_wire3	: STD_LOGIC_VECTOR (31 DOWNTO 0);
	SIGNAL sub_wire4	: STD_LOGIC_VECTOR (31 DOWNTO 0);
	SIGNAL sub_wire5	: STD_LOGIC_VECTOR (31 DOWNTO 0);
	SIGNAL sub_wire6	: STD_LOGIC_VECTOR (31 DOWNTO 0);
	SIGNAL sub_wire7	: STD_LOGIC_VECTOR (31 DOWNTO 0);
	SIGNAL sub_wire8	: STD_LOGIC_VECTOR (31 DOWNTO 0);
	SIGNAL sub_wire9	: STD_LOGIC_VECTOR (31 DOWNTO 0);
	SIGNAL sub_wire10	: STD_LOGIC_VECTOR (31 DOWNTO 0);
	SIGNAL sub_wire11	: STD_LOGIC_VECTOR (31 DOWNTO 0);
	SIGNAL sub_wire12	: STD_LOGIC_VECTOR (31 DOWNTO 0);
	SIGNAL sub_wire13	: STD_LOGIC_VECTOR (31 DOWNTO 0);
	SIGNAL sub_wire14	: STD_LOGIC_VECTOR (31 DOWNTO 0);
	SIGNAL sub_wire15	: STD_LOGIC_VECTOR (31 DOWNTO 0);
	SIGNAL sub_wire16	: STD_LOGIC_VECTOR (31 DOWNTO 0);
	SIGNAL sub_wire17	: STD_LOGIC_VECTOR (31 DOWNTO 0);
	SIGNAL sub_wire18	: STD_LOGIC_VECTOR (31 DOWNTO 0);
	SIGNAL sub_wire19	: STD_LOGIC_VECTOR (31 DOWNTO 0);
	SIGNAL sub_wire20	: STD_LOGIC_VECTOR (31 DOWNTO 0);
	SIGNAL sub_wire21	: STD_LOGIC_VECTOR (31 DOWNTO 0);
	SIGNAL sub_wire22	: STD_LOGIC_VECTOR (31 DOWNTO 0);
	SIGNAL sub_wire23	: STD_LOGIC_VECTOR (31 DOWNTO 0);
	SIGNAL sub_wire24	: STD_LOGIC_VECTOR (31 DOWNTO 0);
	SIGNAL sub_wire25	: STD_LOGIC_VECTOR (31 DOWNTO 0);
	SIGNAL sub_wire26	: STD_LOGIC_VECTOR (31 DOWNTO 0);
	SIGNAL sub_wire27	: STD_LOGIC_VECTOR (31 DOWNTO 0);
	SIGNAL sub_wire28	: STD_LOGIC_VECTOR (31 DOWNTO 0);
	SIGNAL sub_wire29	: STD_LOGIC_VECTOR (31 DOWNTO 0);
	SIGNAL sub_wire30	: STD_LOGIC_VECTOR (31 DOWNTO 0);
	SIGNAL sub_wire31	: STD_LOGIC_VECTOR (31 DOWNTO 0);
	SIGNAL sub_wire32	: STD_LOGIC_VECTOR (31 DOWNTO 0);
	SIGNAL sub_wire33	: STD_LOGIC_VECTOR (31 DOWNTO 0);
	SIGNAL sub_wire34	: STD_LOGIC_VECTOR (31 DOWNTO 0);
	SIGNAL sub_wire35	: STD_LOGIC_VECTOR (31 DOWNTO 0);
	SIGNAL sub_wire36	: STD_LOGIC_VECTOR (31 DOWNTO 0);
	SIGNAL sub_wire37	: STD_LOGIC_VECTOR (31 DOWNTO 0);
	SIGNAL sub_wire38	: STD_LOGIC_VECTOR (31 DOWNTO 0);
	SIGNAL sub_wire39	: STD_LOGIC_VECTOR (31 DOWNTO 0);
	SIGNAL sub_wire40	: STD_LOGIC_VECTOR (31 DOWNTO 0);
	SIGNAL sub_wire41	: STD_LOGIC_VECTOR (31 DOWNTO 0);
	SIGNAL sub_wire42	: STD_LOGIC_VECTOR (31 DOWNTO 0);
	SIGNAL sub_wire43	: STD_LOGIC_VECTOR (31 DOWNTO 0);
	SIGNAL sub_wire44	: STD_LOGIC_VECTOR (31 DOWNTO 0);
	SIGNAL sub_wire45	: STD_LOGIC_VECTOR (31 DOWNTO 0);
	SIGNAL sub_wire46	: STD_LOGIC_VECTOR (31 DOWNTO 0);
	SIGNAL sub_wire47	: STD_LOGIC_VECTOR (31 DOWNTO 0);
	SIGNAL sub_wire48	: STD_LOGIC_VECTOR (31 DOWNTO 0);
	SIGNAL sub_wire49	: STD_LOGIC_VECTOR (31 DOWNTO 0);
	SIGNAL sub_wire50	: STD_LOGIC_VECTOR (31 DOWNTO 0);
	SIGNAL sub_wire51	: STD_LOGIC_VECTOR (31 DOWNTO 0);
	SIGNAL sub_wire52	: STD_LOGIC_VECTOR (31 DOWNTO 0);
	SIGNAL sub_wire53	: STD_LOGIC_VECTOR (31 DOWNTO 0);
	SIGNAL sub_wire54	: STD_LOGIC_VECTOR (31 DOWNTO 0);
	SIGNAL sub_wire55	: STD_LOGIC_VECTOR (31 DOWNTO 0);
	SIGNAL sub_wire56	: STD_LOGIC_VECTOR (31 DOWNTO 0);
	SIGNAL sub_wire57	: STD_LOGIC_VECTOR (31 DOWNTO 0);
	SIGNAL sub_wire58	: STD_LOGIC_VECTOR (31 DOWNTO 0);
	SIGNAL sub_wire59	: STD_LOGIC_VECTOR (31 DOWNTO 0);
	SIGNAL sub_wire60	: STD_LOGIC_VECTOR (31 DOWNTO 0);
	SIGNAL sub_wire61	: STD_LOGIC_VECTOR (31 DOWNTO 0);
	SIGNAL sub_wire62	: STD_LOGIC_VECTOR (31 DOWNTO 0);
	SIGNAL sub_wire63	: STD_LOGIC_VECTOR (31 DOWNTO 0);
	SIGNAL sub_wire64	: STD_LOGIC_VECTOR (31 DOWNTO 0);
	SIGNAL sub_wire65	: STD_LOGIC_VECTOR (31 DOWNTO 0);
	SIGNAL sub_wire66	: STD_LOGIC_VECTOR (31 DOWNTO 0);
	SIGNAL sub_wire67	: STD_LOGIC_VECTOR (31 DOWNTO 0);
	SIGNAL sub_wire68	: STD_LOGIC_VECTOR (31 DOWNTO 0);
	SIGNAL sub_wire69	: STD_LOGIC_VECTOR (31 DOWNTO 0);
	SIGNAL sub_wire70	: STD_LOGIC_VECTOR (31 DOWNTO 0);
	SIGNAL sub_wire71	: STD_LOGIC_VECTOR (31 DOWNTO 0);
	SIGNAL sub_wire72	: STD_LOGIC_VECTOR (31 DOWNTO 0);
	SIGNAL sub_wire73	: STD_LOGIC_VECTOR (31 DOWNTO 0);
	SIGNAL sub_wire74	: STD_LOGIC_VECTOR (31 DOWNTO 0);
	SIGNAL sub_wire75	: STD_LOGIC_VECTOR (31 DOWNTO 0);
	SIGNAL sub_wire76	: STD_LOGIC_VECTOR (31 DOWNTO 0);
	SIGNAL sub_wire77	: STD_LOGIC_VECTOR (31 DOWNTO 0);
	SIGNAL sub_wire78	: STD_LOGIC_VECTOR (31 DOWNTO 0);
	SIGNAL sub_wire79	: STD_LOGIC_VECTOR (31 DOWNTO 0);
	SIGNAL sub_wire80	: STD_LOGIC_VECTOR (31 DOWNTO 0);
	SIGNAL sub_wire81	: STD_LOGIC_VECTOR (31 DOWNTO 0);
	SIGNAL sub_wire82	: STD_LOGIC_VECTOR (31 DOWNTO 0);
	SIGNAL sub_wire83	: STD_LOGIC_VECTOR (31 DOWNTO 0);
	SIGNAL sub_wire84	: STD_LOGIC_VECTOR (31 DOWNTO 0);
	SIGNAL sub_wire85	: STD_LOGIC_VECTOR (31 DOWNTO 0);
	SIGNAL sub_wire86	: STD_LOGIC_VECTOR (31 DOWNTO 0);
	SIGNAL sub_wire87	: STD_LOGIC_VECTOR (31 DOWNTO 0);
	SIGNAL sub_wire88	: STD_LOGIC_VECTOR (31 DOWNTO 0);
	SIGNAL sub_wire89	: STD_LOGIC_VECTOR (31 DOWNTO 0);
	SIGNAL sub_wire90	: STD_LOGIC_VECTOR (31 DOWNTO 0);
	SIGNAL sub_wire91	: STD_LOGIC_VECTOR (31 DOWNTO 0);
	SIGNAL sub_wire92	: STD_LOGIC_VECTOR (31 DOWNTO 0);
	SIGNAL sub_wire93	: STD_LOGIC_VECTOR (31 DOWNTO 0);
	SIGNAL sub_wire94	: STD_LOGIC_VECTOR (31 DOWNTO 0);
	SIGNAL sub_wire95	: STD_LOGIC_VECTOR (31 DOWNTO 0);
	SIGNAL sub_wire96	: STD_LOGIC_VECTOR (31 DOWNTO 0);
	SIGNAL sub_wire97	: STD_LOGIC_VECTOR (31 DOWNTO 0);
	SIGNAL sub_wire98	: STD_LOGIC_VECTOR (31 DOWNTO 0);
	SIGNAL sub_wire99	: STD_LOGIC_VECTOR (31 DOWNTO 0);
	SIGNAL sub_wire100	: STD_LOGIC_VECTOR (31 DOWNTO 0);
	SIGNAL sub_wire101	: STD_LOGIC_VECTOR (31 DOWNTO 0);
	SIGNAL sub_wire102	: STD_LOGIC_VECTOR (31 DOWNTO 0);
	SIGNAL sub_wire103	: STD_LOGIC_VECTOR (31 DOWNTO 0);
	SIGNAL sub_wire104	: STD_LOGIC_VECTOR (31 DOWNTO 0);
	SIGNAL sub_wire105	: STD_LOGIC_VECTOR (31 DOWNTO 0);
	SIGNAL sub_wire106	: STD_LOGIC_VECTOR (31 DOWNTO 0);
	SIGNAL sub_wire107	: STD_LOGIC_VECTOR (31 DOWNTO 0);
	SIGNAL sub_wire108	: STD_LOGIC_VECTOR (31 DOWNTO 0);
	SIGNAL sub_wire109	: STD_LOGIC_VECTOR (31 DOWNTO 0);
	SIGNAL sub_wire110	: STD_LOGIC_VECTOR (31 DOWNTO 0);
	SIGNAL sub_wire111	: STD_LOGIC_VECTOR (31 DOWNTO 0);
	SIGNAL sub_wire112	: STD_LOGIC_VECTOR (31 DOWNTO 0);
	SIGNAL sub_wire113	: STD_LOGIC_VECTOR (31 DOWNTO 0);
	SIGNAL sub_wire114	: STD_LOGIC_VECTOR (31 DOWNTO 0);
	SIGNAL sub_wire115	: STD_LOGIC_VECTOR (31 DOWNTO 0);
	SIGNAL sub_wire116	: STD_LOGIC_VECTOR (31 DOWNTO 0);
	SIGNAL sub_wire117	: STD_LOGIC_VECTOR (31 DOWNTO 0);
	SIGNAL sub_wire118	: STD_LOGIC_VECTOR (31 DOWNTO 0);
	SIGNAL sub_wire119	: STD_LOGIC_VECTOR (31 DOWNTO 0);
	SIGNAL sub_wire120	: STD_LOGIC_VECTOR (31 DOWNTO 0);
	SIGNAL sub_wire121	: STD_LOGIC_VECTOR (31 DOWNTO 0);
	SIGNAL sub_wire122	: STD_LOGIC_VECTOR (31 DOWNTO 0);
	SIGNAL sub_wire123	: STD_LOGIC_VECTOR (31 DOWNTO 0);
	SIGNAL sub_wire124	: STD_LOGIC_VECTOR (31 DOWNTO 0);
	SIGNAL sub_wire125	: STD_LOGIC_VECTOR (31 DOWNTO 0);
	SIGNAL sub_wire126	: STD_LOGIC_VECTOR (31 DOWNTO 0);
	SIGNAL sub_wire127	: STD_LOGIC_VECTOR (31 DOWNTO 0);
	SIGNAL sub_wire128	: STD_LOGIC_VECTOR (31 DOWNTO 0);
	SIGNAL sub_wire129	: STD_LOGIC_VECTOR (31 DOWNTO 0);

BEGIN
	sub_wire128    <= data0x(31 DOWNTO 0);
	sub_wire127    <= data1x(31 DOWNTO 0);
	sub_wire126    <= data2x(31 DOWNTO 0);
	sub_wire125    <= data3x(31 DOWNTO 0);
	sub_wire124    <= data4x(31 DOWNTO 0);
	sub_wire123    <= data5x(31 DOWNTO 0);
	sub_wire122    <= data6x(31 DOWNTO 0);
	sub_wire121    <= data7x(31 DOWNTO 0);
	sub_wire120    <= data8x(31 DOWNTO 0);
	sub_wire119    <= data9x(31 DOWNTO 0);
	sub_wire118    <= data10x(31 DOWNTO 0);
	sub_wire117    <= data11x(31 DOWNTO 0);
	sub_wire116    <= data12x(31 DOWNTO 0);
	sub_wire115    <= data13x(31 DOWNTO 0);
	sub_wire114    <= data14x(31 DOWNTO 0);
	sub_wire113    <= data15x(31 DOWNTO 0);
	sub_wire112    <= data16x(31 DOWNTO 0);
	sub_wire111    <= data17x(31 DOWNTO 0);
	sub_wire110    <= data18x(31 DOWNTO 0);
	sub_wire109    <= data19x(31 DOWNTO 0);
	sub_wire108    <= data20x(31 DOWNTO 0);
	sub_wire107    <= data21x(31 DOWNTO 0);
	sub_wire106    <= data22x(31 DOWNTO 0);
	sub_wire105    <= data23x(31 DOWNTO 0);
	sub_wire104    <= data24x(31 DOWNTO 0);
	sub_wire103    <= data25x(31 DOWNTO 0);
	sub_wire102    <= data26x(31 DOWNTO 0);
	sub_wire101    <= data27x(31 DOWNTO 0);
	sub_wire100    <= data28x(31 DOWNTO 0);
	sub_wire99    <= data29x(31 DOWNTO 0);
	sub_wire98    <= data30x(31 DOWNTO 0);
	sub_wire97    <= data31x(31 DOWNTO 0);
	sub_wire96    <= data32x(31 DOWNTO 0);
	sub_wire95    <= data33x(31 DOWNTO 0);
	sub_wire94    <= data34x(31 DOWNTO 0);
	sub_wire93    <= data35x(31 DOWNTO 0);
	sub_wire92    <= data36x(31 DOWNTO 0);
	sub_wire91    <= data37x(31 DOWNTO 0);
	sub_wire90    <= data38x(31 DOWNTO 0);
	sub_wire89    <= data39x(31 DOWNTO 0);
	sub_wire88    <= data40x(31 DOWNTO 0);
	sub_wire87    <= data41x(31 DOWNTO 0);
	sub_wire86    <= data42x(31 DOWNTO 0);
	sub_wire85    <= data43x(31 DOWNTO 0);
	sub_wire84    <= data44x(31 DOWNTO 0);
	sub_wire83    <= data45x(31 DOWNTO 0);
	sub_wire82    <= data46x(31 DOWNTO 0);
	sub_wire81    <= data47x(31 DOWNTO 0);
	sub_wire80    <= data48x(31 DOWNTO 0);
	sub_wire79    <= data49x(31 DOWNTO 0);
	sub_wire78    <= data50x(31 DOWNTO 0);
	sub_wire77    <= data51x(31 DOWNTO 0);
	sub_wire76    <= data52x(31 DOWNTO 0);
	sub_wire75    <= data53x(31 DOWNTO 0);
	sub_wire74    <= data54x(31 DOWNTO 0);
	sub_wire73    <= data55x(31 DOWNTO 0);
	sub_wire72    <= data56x(31 DOWNTO 0);
	sub_wire71    <= data57x(31 DOWNTO 0);
	sub_wire70    <= data58x(31 DOWNTO 0);
	sub_wire69    <= data59x(31 DOWNTO 0);
	sub_wire68    <= data60x(31 DOWNTO 0);
	sub_wire67    <= data61x(31 DOWNTO 0);
	sub_wire66    <= data62x(31 DOWNTO 0);
	sub_wire65    <= data63x(31 DOWNTO 0);
	sub_wire64    <= data64x(31 DOWNTO 0);
	sub_wire63    <= data65x(31 DOWNTO 0);
	sub_wire62    <= data66x(31 DOWNTO 0);
	sub_wire61    <= data67x(31 DOWNTO 0);
	sub_wire60    <= data68x(31 DOWNTO 0);
	sub_wire59    <= data69x(31 DOWNTO 0);
	sub_wire58    <= data70x(31 DOWNTO 0);
	sub_wire57    <= data71x(31 DOWNTO 0);
	sub_wire56    <= data72x(31 DOWNTO 0);
	sub_wire55    <= data73x(31 DOWNTO 0);
	sub_wire54    <= data74x(31 DOWNTO 0);
	sub_wire53    <= data75x(31 DOWNTO 0);
	sub_wire52    <= data76x(31 DOWNTO 0);
	sub_wire51    <= data77x(31 DOWNTO 0);
	sub_wire50    <= data78x(31 DOWNTO 0);
	sub_wire49    <= data79x(31 DOWNTO 0);
	sub_wire48    <= data80x(31 DOWNTO 0);
	sub_wire47    <= data81x(31 DOWNTO 0);
	sub_wire46    <= data82x(31 DOWNTO 0);
	sub_wire45    <= data83x(31 DOWNTO 0);
	sub_wire44    <= data84x(31 DOWNTO 0);
	sub_wire43    <= data85x(31 DOWNTO 0);
	sub_wire42    <= data86x(31 DOWNTO 0);
	sub_wire41    <= data87x(31 DOWNTO 0);
	sub_wire40    <= data88x(31 DOWNTO 0);
	sub_wire39    <= data89x(31 DOWNTO 0);
	sub_wire38    <= data90x(31 DOWNTO 0);
	sub_wire37    <= data91x(31 DOWNTO 0);
	sub_wire36    <= data92x(31 DOWNTO 0);
	sub_wire35    <= data93x(31 DOWNTO 0);
	sub_wire34    <= data94x(31 DOWNTO 0);
	sub_wire33    <= data95x(31 DOWNTO 0);
	sub_wire32    <= data96x(31 DOWNTO 0);
	sub_wire31    <= data97x(31 DOWNTO 0);
	sub_wire30    <= data98x(31 DOWNTO 0);
	sub_wire29    <= data99x(31 DOWNTO 0);
	sub_wire28    <= data100x(31 DOWNTO 0);
	sub_wire27    <= data101x(31 DOWNTO 0);
	sub_wire26    <= data102x(31 DOWNTO 0);
	sub_wire25    <= data103x(31 DOWNTO 0);
	sub_wire24    <= data104x(31 DOWNTO 0);
	sub_wire23    <= data105x(31 DOWNTO 0);
	sub_wire22    <= data106x(31 DOWNTO 0);
	sub_wire21    <= data107x(31 DOWNTO 0);
	sub_wire20    <= data108x(31 DOWNTO 0);
	sub_wire19    <= data109x(31 DOWNTO 0);
	sub_wire18    <= data110x(31 DOWNTO 0);
	sub_wire17    <= data111x(31 DOWNTO 0);
	sub_wire16    <= data112x(31 DOWNTO 0);
	sub_wire15    <= data113x(31 DOWNTO 0);
	sub_wire14    <= data114x(31 DOWNTO 0);
	sub_wire13    <= data115x(31 DOWNTO 0);
	sub_wire12    <= data116x(31 DOWNTO 0);
	sub_wire11    <= data117x(31 DOWNTO 0);
	sub_wire10    <= data118x(31 DOWNTO 0);
	sub_wire9    <= data119x(31 DOWNTO 0);
	sub_wire8    <= data120x(31 DOWNTO 0);
	sub_wire7    <= data121x(31 DOWNTO 0);
	sub_wire6    <= data122x(31 DOWNTO 0);
	sub_wire5    <= data123x(31 DOWNTO 0);
	sub_wire4    <= data124x(31 DOWNTO 0);
	sub_wire3    <= data125x(31 DOWNTO 0);
	sub_wire2    <= data126x(31 DOWNTO 0);
	sub_wire0    <= data127x(31 DOWNTO 0);
	sub_wire1(127, 0)    <= sub_wire0(0);
	sub_wire1(127, 1)    <= sub_wire0(1);
	sub_wire1(127, 2)    <= sub_wire0(2);
	sub_wire1(127, 3)    <= sub_wire0(3);
	sub_wire1(127, 4)    <= sub_wire0(4);
	sub_wire1(127, 5)    <= sub_wire0(5);
	sub_wire1(127, 6)    <= sub_wire0(6);
	sub_wire1(127, 7)    <= sub_wire0(7);
	sub_wire1(127, 8)    <= sub_wire0(8);
	sub_wire1(127, 9)    <= sub_wire0(9);
	sub_wire1(127, 10)    <= sub_wire0(10);
	sub_wire1(127, 11)    <= sub_wire0(11);
	sub_wire1(127, 12)    <= sub_wire0(12);
	sub_wire1(127, 13)    <= sub_wire0(13);
	sub_wire1(127, 14)    <= sub_wire0(14);
	sub_wire1(127, 15)    <= sub_wire0(15);
	sub_wire1(127, 16)    <= sub_wire0(16);
	sub_wire1(127, 17)    <= sub_wire0(17);
	sub_wire1(127, 18)    <= sub_wire0(18);
	sub_wire1(127, 19)    <= sub_wire0(19);
	sub_wire1(127, 20)    <= sub_wire0(20);
	sub_wire1(127, 21)    <= sub_wire0(21);
	sub_wire1(127, 22)    <= sub_wire0(22);
	sub_wire1(127, 23)    <= sub_wire0(23);
	sub_wire1(127, 24)    <= sub_wire0(24);
	sub_wire1(127, 25)    <= sub_wire0(25);
	sub_wire1(127, 26)    <= sub_wire0(26);
	sub_wire1(127, 27)    <= sub_wire0(27);
	sub_wire1(127, 28)    <= sub_wire0(28);
	sub_wire1(127, 29)    <= sub_wire0(29);
	sub_wire1(127, 30)    <= sub_wire0(30);
	sub_wire1(127, 31)    <= sub_wire0(31);
	sub_wire1(126, 0)    <= sub_wire2(0);
	sub_wire1(126, 1)    <= sub_wire2(1);
	sub_wire1(126, 2)    <= sub_wire2(2);
	sub_wire1(126, 3)    <= sub_wire2(3);
	sub_wire1(126, 4)    <= sub_wire2(4);
	sub_wire1(126, 5)    <= sub_wire2(5);
	sub_wire1(126, 6)    <= sub_wire2(6);
	sub_wire1(126, 7)    <= sub_wire2(7);
	sub_wire1(126, 8)    <= sub_wire2(8);
	sub_wire1(126, 9)    <= sub_wire2(9);
	sub_wire1(126, 10)    <= sub_wire2(10);
	sub_wire1(126, 11)    <= sub_wire2(11);
	sub_wire1(126, 12)    <= sub_wire2(12);
	sub_wire1(126, 13)    <= sub_wire2(13);
	sub_wire1(126, 14)    <= sub_wire2(14);
	sub_wire1(126, 15)    <= sub_wire2(15);
	sub_wire1(126, 16)    <= sub_wire2(16);
	sub_wire1(126, 17)    <= sub_wire2(17);
	sub_wire1(126, 18)    <= sub_wire2(18);
	sub_wire1(126, 19)    <= sub_wire2(19);
	sub_wire1(126, 20)    <= sub_wire2(20);
	sub_wire1(126, 21)    <= sub_wire2(21);
	sub_wire1(126, 22)    <= sub_wire2(22);
	sub_wire1(126, 23)    <= sub_wire2(23);
	sub_wire1(126, 24)    <= sub_wire2(24);
	sub_wire1(126, 25)    <= sub_wire2(25);
	sub_wire1(126, 26)    <= sub_wire2(26);
	sub_wire1(126, 27)    <= sub_wire2(27);
	sub_wire1(126, 28)    <= sub_wire2(28);
	sub_wire1(126, 29)    <= sub_wire2(29);
	sub_wire1(126, 30)    <= sub_wire2(30);
	sub_wire1(126, 31)    <= sub_wire2(31);
	sub_wire1(125, 0)    <= sub_wire3(0);
	sub_wire1(125, 1)    <= sub_wire3(1);
	sub_wire1(125, 2)    <= sub_wire3(2);
	sub_wire1(125, 3)    <= sub_wire3(3);
	sub_wire1(125, 4)    <= sub_wire3(4);
	sub_wire1(125, 5)    <= sub_wire3(5);
	sub_wire1(125, 6)    <= sub_wire3(6);
	sub_wire1(125, 7)    <= sub_wire3(7);
	sub_wire1(125, 8)    <= sub_wire3(8);
	sub_wire1(125, 9)    <= sub_wire3(9);
	sub_wire1(125, 10)    <= sub_wire3(10);
	sub_wire1(125, 11)    <= sub_wire3(11);
	sub_wire1(125, 12)    <= sub_wire3(12);
	sub_wire1(125, 13)    <= sub_wire3(13);
	sub_wire1(125, 14)    <= sub_wire3(14);
	sub_wire1(125, 15)    <= sub_wire3(15);
	sub_wire1(125, 16)    <= sub_wire3(16);
	sub_wire1(125, 17)    <= sub_wire3(17);
	sub_wire1(125, 18)    <= sub_wire3(18);
	sub_wire1(125, 19)    <= sub_wire3(19);
	sub_wire1(125, 20)    <= sub_wire3(20);
	sub_wire1(125, 21)    <= sub_wire3(21);
	sub_wire1(125, 22)    <= sub_wire3(22);
	sub_wire1(125, 23)    <= sub_wire3(23);
	sub_wire1(125, 24)    <= sub_wire3(24);
	sub_wire1(125, 25)    <= sub_wire3(25);
	sub_wire1(125, 26)    <= sub_wire3(26);
	sub_wire1(125, 27)    <= sub_wire3(27);
	sub_wire1(125, 28)    <= sub_wire3(28);
	sub_wire1(125, 29)    <= sub_wire3(29);
	sub_wire1(125, 30)    <= sub_wire3(30);
	sub_wire1(125, 31)    <= sub_wire3(31);
	sub_wire1(124, 0)    <= sub_wire4(0);
	sub_wire1(124, 1)    <= sub_wire4(1);
	sub_wire1(124, 2)    <= sub_wire4(2);
	sub_wire1(124, 3)    <= sub_wire4(3);
	sub_wire1(124, 4)    <= sub_wire4(4);
	sub_wire1(124, 5)    <= sub_wire4(5);
	sub_wire1(124, 6)    <= sub_wire4(6);
	sub_wire1(124, 7)    <= sub_wire4(7);
	sub_wire1(124, 8)    <= sub_wire4(8);
	sub_wire1(124, 9)    <= sub_wire4(9);
	sub_wire1(124, 10)    <= sub_wire4(10);
	sub_wire1(124, 11)    <= sub_wire4(11);
	sub_wire1(124, 12)    <= sub_wire4(12);
	sub_wire1(124, 13)    <= sub_wire4(13);
	sub_wire1(124, 14)    <= sub_wire4(14);
	sub_wire1(124, 15)    <= sub_wire4(15);
	sub_wire1(124, 16)    <= sub_wire4(16);
	sub_wire1(124, 17)    <= sub_wire4(17);
	sub_wire1(124, 18)    <= sub_wire4(18);
	sub_wire1(124, 19)    <= sub_wire4(19);
	sub_wire1(124, 20)    <= sub_wire4(20);
	sub_wire1(124, 21)    <= sub_wire4(21);
	sub_wire1(124, 22)    <= sub_wire4(22);
	sub_wire1(124, 23)    <= sub_wire4(23);
	sub_wire1(124, 24)    <= sub_wire4(24);
	sub_wire1(124, 25)    <= sub_wire4(25);
	sub_wire1(124, 26)    <= sub_wire4(26);
	sub_wire1(124, 27)    <= sub_wire4(27);
	sub_wire1(124, 28)    <= sub_wire4(28);
	sub_wire1(124, 29)    <= sub_wire4(29);
	sub_wire1(124, 30)    <= sub_wire4(30);
	sub_wire1(124, 31)    <= sub_wire4(31);
	sub_wire1(123, 0)    <= sub_wire5(0);
	sub_wire1(123, 1)    <= sub_wire5(1);
	sub_wire1(123, 2)    <= sub_wire5(2);
	sub_wire1(123, 3)    <= sub_wire5(3);
	sub_wire1(123, 4)    <= sub_wire5(4);
	sub_wire1(123, 5)    <= sub_wire5(5);
	sub_wire1(123, 6)    <= sub_wire5(6);
	sub_wire1(123, 7)    <= sub_wire5(7);
	sub_wire1(123, 8)    <= sub_wire5(8);
	sub_wire1(123, 9)    <= sub_wire5(9);
	sub_wire1(123, 10)    <= sub_wire5(10);
	sub_wire1(123, 11)    <= sub_wire5(11);
	sub_wire1(123, 12)    <= sub_wire5(12);
	sub_wire1(123, 13)    <= sub_wire5(13);
	sub_wire1(123, 14)    <= sub_wire5(14);
	sub_wire1(123, 15)    <= sub_wire5(15);
	sub_wire1(123, 16)    <= sub_wire5(16);
	sub_wire1(123, 17)    <= sub_wire5(17);
	sub_wire1(123, 18)    <= sub_wire5(18);
	sub_wire1(123, 19)    <= sub_wire5(19);
	sub_wire1(123, 20)    <= sub_wire5(20);
	sub_wire1(123, 21)    <= sub_wire5(21);
	sub_wire1(123, 22)    <= sub_wire5(22);
	sub_wire1(123, 23)    <= sub_wire5(23);
	sub_wire1(123, 24)    <= sub_wire5(24);
	sub_wire1(123, 25)    <= sub_wire5(25);
	sub_wire1(123, 26)    <= sub_wire5(26);
	sub_wire1(123, 27)    <= sub_wire5(27);
	sub_wire1(123, 28)    <= sub_wire5(28);
	sub_wire1(123, 29)    <= sub_wire5(29);
	sub_wire1(123, 30)    <= sub_wire5(30);
	sub_wire1(123, 31)    <= sub_wire5(31);
	sub_wire1(122, 0)    <= sub_wire6(0);
	sub_wire1(122, 1)    <= sub_wire6(1);
	sub_wire1(122, 2)    <= sub_wire6(2);
	sub_wire1(122, 3)    <= sub_wire6(3);
	sub_wire1(122, 4)    <= sub_wire6(4);
	sub_wire1(122, 5)    <= sub_wire6(5);
	sub_wire1(122, 6)    <= sub_wire6(6);
	sub_wire1(122, 7)    <= sub_wire6(7);
	sub_wire1(122, 8)    <= sub_wire6(8);
	sub_wire1(122, 9)    <= sub_wire6(9);
	sub_wire1(122, 10)    <= sub_wire6(10);
	sub_wire1(122, 11)    <= sub_wire6(11);
	sub_wire1(122, 12)    <= sub_wire6(12);
	sub_wire1(122, 13)    <= sub_wire6(13);
	sub_wire1(122, 14)    <= sub_wire6(14);
	sub_wire1(122, 15)    <= sub_wire6(15);
	sub_wire1(122, 16)    <= sub_wire6(16);
	sub_wire1(122, 17)    <= sub_wire6(17);
	sub_wire1(122, 18)    <= sub_wire6(18);
	sub_wire1(122, 19)    <= sub_wire6(19);
	sub_wire1(122, 20)    <= sub_wire6(20);
	sub_wire1(122, 21)    <= sub_wire6(21);
	sub_wire1(122, 22)    <= sub_wire6(22);
	sub_wire1(122, 23)    <= sub_wire6(23);
	sub_wire1(122, 24)    <= sub_wire6(24);
	sub_wire1(122, 25)    <= sub_wire6(25);
	sub_wire1(122, 26)    <= sub_wire6(26);
	sub_wire1(122, 27)    <= sub_wire6(27);
	sub_wire1(122, 28)    <= sub_wire6(28);
	sub_wire1(122, 29)    <= sub_wire6(29);
	sub_wire1(122, 30)    <= sub_wire6(30);
	sub_wire1(122, 31)    <= sub_wire6(31);
	sub_wire1(121, 0)    <= sub_wire7(0);
	sub_wire1(121, 1)    <= sub_wire7(1);
	sub_wire1(121, 2)    <= sub_wire7(2);
	sub_wire1(121, 3)    <= sub_wire7(3);
	sub_wire1(121, 4)    <= sub_wire7(4);
	sub_wire1(121, 5)    <= sub_wire7(5);
	sub_wire1(121, 6)    <= sub_wire7(6);
	sub_wire1(121, 7)    <= sub_wire7(7);
	sub_wire1(121, 8)    <= sub_wire7(8);
	sub_wire1(121, 9)    <= sub_wire7(9);
	sub_wire1(121, 10)    <= sub_wire7(10);
	sub_wire1(121, 11)    <= sub_wire7(11);
	sub_wire1(121, 12)    <= sub_wire7(12);
	sub_wire1(121, 13)    <= sub_wire7(13);
	sub_wire1(121, 14)    <= sub_wire7(14);
	sub_wire1(121, 15)    <= sub_wire7(15);
	sub_wire1(121, 16)    <= sub_wire7(16);
	sub_wire1(121, 17)    <= sub_wire7(17);
	sub_wire1(121, 18)    <= sub_wire7(18);
	sub_wire1(121, 19)    <= sub_wire7(19);
	sub_wire1(121, 20)    <= sub_wire7(20);
	sub_wire1(121, 21)    <= sub_wire7(21);
	sub_wire1(121, 22)    <= sub_wire7(22);
	sub_wire1(121, 23)    <= sub_wire7(23);
	sub_wire1(121, 24)    <= sub_wire7(24);
	sub_wire1(121, 25)    <= sub_wire7(25);
	sub_wire1(121, 26)    <= sub_wire7(26);
	sub_wire1(121, 27)    <= sub_wire7(27);
	sub_wire1(121, 28)    <= sub_wire7(28);
	sub_wire1(121, 29)    <= sub_wire7(29);
	sub_wire1(121, 30)    <= sub_wire7(30);
	sub_wire1(121, 31)    <= sub_wire7(31);
	sub_wire1(120, 0)    <= sub_wire8(0);
	sub_wire1(120, 1)    <= sub_wire8(1);
	sub_wire1(120, 2)    <= sub_wire8(2);
	sub_wire1(120, 3)    <= sub_wire8(3);
	sub_wire1(120, 4)    <= sub_wire8(4);
	sub_wire1(120, 5)    <= sub_wire8(5);
	sub_wire1(120, 6)    <= sub_wire8(6);
	sub_wire1(120, 7)    <= sub_wire8(7);
	sub_wire1(120, 8)    <= sub_wire8(8);
	sub_wire1(120, 9)    <= sub_wire8(9);
	sub_wire1(120, 10)    <= sub_wire8(10);
	sub_wire1(120, 11)    <= sub_wire8(11);
	sub_wire1(120, 12)    <= sub_wire8(12);
	sub_wire1(120, 13)    <= sub_wire8(13);
	sub_wire1(120, 14)    <= sub_wire8(14);
	sub_wire1(120, 15)    <= sub_wire8(15);
	sub_wire1(120, 16)    <= sub_wire8(16);
	sub_wire1(120, 17)    <= sub_wire8(17);
	sub_wire1(120, 18)    <= sub_wire8(18);
	sub_wire1(120, 19)    <= sub_wire8(19);
	sub_wire1(120, 20)    <= sub_wire8(20);
	sub_wire1(120, 21)    <= sub_wire8(21);
	sub_wire1(120, 22)    <= sub_wire8(22);
	sub_wire1(120, 23)    <= sub_wire8(23);
	sub_wire1(120, 24)    <= sub_wire8(24);
	sub_wire1(120, 25)    <= sub_wire8(25);
	sub_wire1(120, 26)    <= sub_wire8(26);
	sub_wire1(120, 27)    <= sub_wire8(27);
	sub_wire1(120, 28)    <= sub_wire8(28);
	sub_wire1(120, 29)    <= sub_wire8(29);
	sub_wire1(120, 30)    <= sub_wire8(30);
	sub_wire1(120, 31)    <= sub_wire8(31);
	sub_wire1(119, 0)    <= sub_wire9(0);
	sub_wire1(119, 1)    <= sub_wire9(1);
	sub_wire1(119, 2)    <= sub_wire9(2);
	sub_wire1(119, 3)    <= sub_wire9(3);
	sub_wire1(119, 4)    <= sub_wire9(4);
	sub_wire1(119, 5)    <= sub_wire9(5);
	sub_wire1(119, 6)    <= sub_wire9(6);
	sub_wire1(119, 7)    <= sub_wire9(7);
	sub_wire1(119, 8)    <= sub_wire9(8);
	sub_wire1(119, 9)    <= sub_wire9(9);
	sub_wire1(119, 10)    <= sub_wire9(10);
	sub_wire1(119, 11)    <= sub_wire9(11);
	sub_wire1(119, 12)    <= sub_wire9(12);
	sub_wire1(119, 13)    <= sub_wire9(13);
	sub_wire1(119, 14)    <= sub_wire9(14);
	sub_wire1(119, 15)    <= sub_wire9(15);
	sub_wire1(119, 16)    <= sub_wire9(16);
	sub_wire1(119, 17)    <= sub_wire9(17);
	sub_wire1(119, 18)    <= sub_wire9(18);
	sub_wire1(119, 19)    <= sub_wire9(19);
	sub_wire1(119, 20)    <= sub_wire9(20);
	sub_wire1(119, 21)    <= sub_wire9(21);
	sub_wire1(119, 22)    <= sub_wire9(22);
	sub_wire1(119, 23)    <= sub_wire9(23);
	sub_wire1(119, 24)    <= sub_wire9(24);
	sub_wire1(119, 25)    <= sub_wire9(25);
	sub_wire1(119, 26)    <= sub_wire9(26);
	sub_wire1(119, 27)    <= sub_wire9(27);
	sub_wire1(119, 28)    <= sub_wire9(28);
	sub_wire1(119, 29)    <= sub_wire9(29);
	sub_wire1(119, 30)    <= sub_wire9(30);
	sub_wire1(119, 31)    <= sub_wire9(31);
	sub_wire1(118, 0)    <= sub_wire10(0);
	sub_wire1(118, 1)    <= sub_wire10(1);
	sub_wire1(118, 2)    <= sub_wire10(2);
	sub_wire1(118, 3)    <= sub_wire10(3);
	sub_wire1(118, 4)    <= sub_wire10(4);
	sub_wire1(118, 5)    <= sub_wire10(5);
	sub_wire1(118, 6)    <= sub_wire10(6);
	sub_wire1(118, 7)    <= sub_wire10(7);
	sub_wire1(118, 8)    <= sub_wire10(8);
	sub_wire1(118, 9)    <= sub_wire10(9);
	sub_wire1(118, 10)    <= sub_wire10(10);
	sub_wire1(118, 11)    <= sub_wire10(11);
	sub_wire1(118, 12)    <= sub_wire10(12);
	sub_wire1(118, 13)    <= sub_wire10(13);
	sub_wire1(118, 14)    <= sub_wire10(14);
	sub_wire1(118, 15)    <= sub_wire10(15);
	sub_wire1(118, 16)    <= sub_wire10(16);
	sub_wire1(118, 17)    <= sub_wire10(17);
	sub_wire1(118, 18)    <= sub_wire10(18);
	sub_wire1(118, 19)    <= sub_wire10(19);
	sub_wire1(118, 20)    <= sub_wire10(20);
	sub_wire1(118, 21)    <= sub_wire10(21);
	sub_wire1(118, 22)    <= sub_wire10(22);
	sub_wire1(118, 23)    <= sub_wire10(23);
	sub_wire1(118, 24)    <= sub_wire10(24);
	sub_wire1(118, 25)    <= sub_wire10(25);
	sub_wire1(118, 26)    <= sub_wire10(26);
	sub_wire1(118, 27)    <= sub_wire10(27);
	sub_wire1(118, 28)    <= sub_wire10(28);
	sub_wire1(118, 29)    <= sub_wire10(29);
	sub_wire1(118, 30)    <= sub_wire10(30);
	sub_wire1(118, 31)    <= sub_wire10(31);
	sub_wire1(117, 0)    <= sub_wire11(0);
	sub_wire1(117, 1)    <= sub_wire11(1);
	sub_wire1(117, 2)    <= sub_wire11(2);
	sub_wire1(117, 3)    <= sub_wire11(3);
	sub_wire1(117, 4)    <= sub_wire11(4);
	sub_wire1(117, 5)    <= sub_wire11(5);
	sub_wire1(117, 6)    <= sub_wire11(6);
	sub_wire1(117, 7)    <= sub_wire11(7);
	sub_wire1(117, 8)    <= sub_wire11(8);
	sub_wire1(117, 9)    <= sub_wire11(9);
	sub_wire1(117, 10)    <= sub_wire11(10);
	sub_wire1(117, 11)    <= sub_wire11(11);
	sub_wire1(117, 12)    <= sub_wire11(12);
	sub_wire1(117, 13)    <= sub_wire11(13);
	sub_wire1(117, 14)    <= sub_wire11(14);
	sub_wire1(117, 15)    <= sub_wire11(15);
	sub_wire1(117, 16)    <= sub_wire11(16);
	sub_wire1(117, 17)    <= sub_wire11(17);
	sub_wire1(117, 18)    <= sub_wire11(18);
	sub_wire1(117, 19)    <= sub_wire11(19);
	sub_wire1(117, 20)    <= sub_wire11(20);
	sub_wire1(117, 21)    <= sub_wire11(21);
	sub_wire1(117, 22)    <= sub_wire11(22);
	sub_wire1(117, 23)    <= sub_wire11(23);
	sub_wire1(117, 24)    <= sub_wire11(24);
	sub_wire1(117, 25)    <= sub_wire11(25);
	sub_wire1(117, 26)    <= sub_wire11(26);
	sub_wire1(117, 27)    <= sub_wire11(27);
	sub_wire1(117, 28)    <= sub_wire11(28);
	sub_wire1(117, 29)    <= sub_wire11(29);
	sub_wire1(117, 30)    <= sub_wire11(30);
	sub_wire1(117, 31)    <= sub_wire11(31);
	sub_wire1(116, 0)    <= sub_wire12(0);
	sub_wire1(116, 1)    <= sub_wire12(1);
	sub_wire1(116, 2)    <= sub_wire12(2);
	sub_wire1(116, 3)    <= sub_wire12(3);
	sub_wire1(116, 4)    <= sub_wire12(4);
	sub_wire1(116, 5)    <= sub_wire12(5);
	sub_wire1(116, 6)    <= sub_wire12(6);
	sub_wire1(116, 7)    <= sub_wire12(7);
	sub_wire1(116, 8)    <= sub_wire12(8);
	sub_wire1(116, 9)    <= sub_wire12(9);
	sub_wire1(116, 10)    <= sub_wire12(10);
	sub_wire1(116, 11)    <= sub_wire12(11);
	sub_wire1(116, 12)    <= sub_wire12(12);
	sub_wire1(116, 13)    <= sub_wire12(13);
	sub_wire1(116, 14)    <= sub_wire12(14);
	sub_wire1(116, 15)    <= sub_wire12(15);
	sub_wire1(116, 16)    <= sub_wire12(16);
	sub_wire1(116, 17)    <= sub_wire12(17);
	sub_wire1(116, 18)    <= sub_wire12(18);
	sub_wire1(116, 19)    <= sub_wire12(19);
	sub_wire1(116, 20)    <= sub_wire12(20);
	sub_wire1(116, 21)    <= sub_wire12(21);
	sub_wire1(116, 22)    <= sub_wire12(22);
	sub_wire1(116, 23)    <= sub_wire12(23);
	sub_wire1(116, 24)    <= sub_wire12(24);
	sub_wire1(116, 25)    <= sub_wire12(25);
	sub_wire1(116, 26)    <= sub_wire12(26);
	sub_wire1(116, 27)    <= sub_wire12(27);
	sub_wire1(116, 28)    <= sub_wire12(28);
	sub_wire1(116, 29)    <= sub_wire12(29);
	sub_wire1(116, 30)    <= sub_wire12(30);
	sub_wire1(116, 31)    <= sub_wire12(31);
	sub_wire1(115, 0)    <= sub_wire13(0);
	sub_wire1(115, 1)    <= sub_wire13(1);
	sub_wire1(115, 2)    <= sub_wire13(2);
	sub_wire1(115, 3)    <= sub_wire13(3);
	sub_wire1(115, 4)    <= sub_wire13(4);
	sub_wire1(115, 5)    <= sub_wire13(5);
	sub_wire1(115, 6)    <= sub_wire13(6);
	sub_wire1(115, 7)    <= sub_wire13(7);
	sub_wire1(115, 8)    <= sub_wire13(8);
	sub_wire1(115, 9)    <= sub_wire13(9);
	sub_wire1(115, 10)    <= sub_wire13(10);
	sub_wire1(115, 11)    <= sub_wire13(11);
	sub_wire1(115, 12)    <= sub_wire13(12);
	sub_wire1(115, 13)    <= sub_wire13(13);
	sub_wire1(115, 14)    <= sub_wire13(14);
	sub_wire1(115, 15)    <= sub_wire13(15);
	sub_wire1(115, 16)    <= sub_wire13(16);
	sub_wire1(115, 17)    <= sub_wire13(17);
	sub_wire1(115, 18)    <= sub_wire13(18);
	sub_wire1(115, 19)    <= sub_wire13(19);
	sub_wire1(115, 20)    <= sub_wire13(20);
	sub_wire1(115, 21)    <= sub_wire13(21);
	sub_wire1(115, 22)    <= sub_wire13(22);
	sub_wire1(115, 23)    <= sub_wire13(23);
	sub_wire1(115, 24)    <= sub_wire13(24);
	sub_wire1(115, 25)    <= sub_wire13(25);
	sub_wire1(115, 26)    <= sub_wire13(26);
	sub_wire1(115, 27)    <= sub_wire13(27);
	sub_wire1(115, 28)    <= sub_wire13(28);
	sub_wire1(115, 29)    <= sub_wire13(29);
	sub_wire1(115, 30)    <= sub_wire13(30);
	sub_wire1(115, 31)    <= sub_wire13(31);
	sub_wire1(114, 0)    <= sub_wire14(0);
	sub_wire1(114, 1)    <= sub_wire14(1);
	sub_wire1(114, 2)    <= sub_wire14(2);
	sub_wire1(114, 3)    <= sub_wire14(3);
	sub_wire1(114, 4)    <= sub_wire14(4);
	sub_wire1(114, 5)    <= sub_wire14(5);
	sub_wire1(114, 6)    <= sub_wire14(6);
	sub_wire1(114, 7)    <= sub_wire14(7);
	sub_wire1(114, 8)    <= sub_wire14(8);
	sub_wire1(114, 9)    <= sub_wire14(9);
	sub_wire1(114, 10)    <= sub_wire14(10);
	sub_wire1(114, 11)    <= sub_wire14(11);
	sub_wire1(114, 12)    <= sub_wire14(12);
	sub_wire1(114, 13)    <= sub_wire14(13);
	sub_wire1(114, 14)    <= sub_wire14(14);
	sub_wire1(114, 15)    <= sub_wire14(15);
	sub_wire1(114, 16)    <= sub_wire14(16);
	sub_wire1(114, 17)    <= sub_wire14(17);
	sub_wire1(114, 18)    <= sub_wire14(18);
	sub_wire1(114, 19)    <= sub_wire14(19);
	sub_wire1(114, 20)    <= sub_wire14(20);
	sub_wire1(114, 21)    <= sub_wire14(21);
	sub_wire1(114, 22)    <= sub_wire14(22);
	sub_wire1(114, 23)    <= sub_wire14(23);
	sub_wire1(114, 24)    <= sub_wire14(24);
	sub_wire1(114, 25)    <= sub_wire14(25);
	sub_wire1(114, 26)    <= sub_wire14(26);
	sub_wire1(114, 27)    <= sub_wire14(27);
	sub_wire1(114, 28)    <= sub_wire14(28);
	sub_wire1(114, 29)    <= sub_wire14(29);
	sub_wire1(114, 30)    <= sub_wire14(30);
	sub_wire1(114, 31)    <= sub_wire14(31);
	sub_wire1(113, 0)    <= sub_wire15(0);
	sub_wire1(113, 1)    <= sub_wire15(1);
	sub_wire1(113, 2)    <= sub_wire15(2);
	sub_wire1(113, 3)    <= sub_wire15(3);
	sub_wire1(113, 4)    <= sub_wire15(4);
	sub_wire1(113, 5)    <= sub_wire15(5);
	sub_wire1(113, 6)    <= sub_wire15(6);
	sub_wire1(113, 7)    <= sub_wire15(7);
	sub_wire1(113, 8)    <= sub_wire15(8);
	sub_wire1(113, 9)    <= sub_wire15(9);
	sub_wire1(113, 10)    <= sub_wire15(10);
	sub_wire1(113, 11)    <= sub_wire15(11);
	sub_wire1(113, 12)    <= sub_wire15(12);
	sub_wire1(113, 13)    <= sub_wire15(13);
	sub_wire1(113, 14)    <= sub_wire15(14);
	sub_wire1(113, 15)    <= sub_wire15(15);
	sub_wire1(113, 16)    <= sub_wire15(16);
	sub_wire1(113, 17)    <= sub_wire15(17);
	sub_wire1(113, 18)    <= sub_wire15(18);
	sub_wire1(113, 19)    <= sub_wire15(19);
	sub_wire1(113, 20)    <= sub_wire15(20);
	sub_wire1(113, 21)    <= sub_wire15(21);
	sub_wire1(113, 22)    <= sub_wire15(22);
	sub_wire1(113, 23)    <= sub_wire15(23);
	sub_wire1(113, 24)    <= sub_wire15(24);
	sub_wire1(113, 25)    <= sub_wire15(25);
	sub_wire1(113, 26)    <= sub_wire15(26);
	sub_wire1(113, 27)    <= sub_wire15(27);
	sub_wire1(113, 28)    <= sub_wire15(28);
	sub_wire1(113, 29)    <= sub_wire15(29);
	sub_wire1(113, 30)    <= sub_wire15(30);
	sub_wire1(113, 31)    <= sub_wire15(31);
	sub_wire1(112, 0)    <= sub_wire16(0);
	sub_wire1(112, 1)    <= sub_wire16(1);
	sub_wire1(112, 2)    <= sub_wire16(2);
	sub_wire1(112, 3)    <= sub_wire16(3);
	sub_wire1(112, 4)    <= sub_wire16(4);
	sub_wire1(112, 5)    <= sub_wire16(5);
	sub_wire1(112, 6)    <= sub_wire16(6);
	sub_wire1(112, 7)    <= sub_wire16(7);
	sub_wire1(112, 8)    <= sub_wire16(8);
	sub_wire1(112, 9)    <= sub_wire16(9);
	sub_wire1(112, 10)    <= sub_wire16(10);
	sub_wire1(112, 11)    <= sub_wire16(11);
	sub_wire1(112, 12)    <= sub_wire16(12);
	sub_wire1(112, 13)    <= sub_wire16(13);
	sub_wire1(112, 14)    <= sub_wire16(14);
	sub_wire1(112, 15)    <= sub_wire16(15);
	sub_wire1(112, 16)    <= sub_wire16(16);
	sub_wire1(112, 17)    <= sub_wire16(17);
	sub_wire1(112, 18)    <= sub_wire16(18);
	sub_wire1(112, 19)    <= sub_wire16(19);
	sub_wire1(112, 20)    <= sub_wire16(20);
	sub_wire1(112, 21)    <= sub_wire16(21);
	sub_wire1(112, 22)    <= sub_wire16(22);
	sub_wire1(112, 23)    <= sub_wire16(23);
	sub_wire1(112, 24)    <= sub_wire16(24);
	sub_wire1(112, 25)    <= sub_wire16(25);
	sub_wire1(112, 26)    <= sub_wire16(26);
	sub_wire1(112, 27)    <= sub_wire16(27);
	sub_wire1(112, 28)    <= sub_wire16(28);
	sub_wire1(112, 29)    <= sub_wire16(29);
	sub_wire1(112, 30)    <= sub_wire16(30);
	sub_wire1(112, 31)    <= sub_wire16(31);
	sub_wire1(111, 0)    <= sub_wire17(0);
	sub_wire1(111, 1)    <= sub_wire17(1);
	sub_wire1(111, 2)    <= sub_wire17(2);
	sub_wire1(111, 3)    <= sub_wire17(3);
	sub_wire1(111, 4)    <= sub_wire17(4);
	sub_wire1(111, 5)    <= sub_wire17(5);
	sub_wire1(111, 6)    <= sub_wire17(6);
	sub_wire1(111, 7)    <= sub_wire17(7);
	sub_wire1(111, 8)    <= sub_wire17(8);
	sub_wire1(111, 9)    <= sub_wire17(9);
	sub_wire1(111, 10)    <= sub_wire17(10);
	sub_wire1(111, 11)    <= sub_wire17(11);
	sub_wire1(111, 12)    <= sub_wire17(12);
	sub_wire1(111, 13)    <= sub_wire17(13);
	sub_wire1(111, 14)    <= sub_wire17(14);
	sub_wire1(111, 15)    <= sub_wire17(15);
	sub_wire1(111, 16)    <= sub_wire17(16);
	sub_wire1(111, 17)    <= sub_wire17(17);
	sub_wire1(111, 18)    <= sub_wire17(18);
	sub_wire1(111, 19)    <= sub_wire17(19);
	sub_wire1(111, 20)    <= sub_wire17(20);
	sub_wire1(111, 21)    <= sub_wire17(21);
	sub_wire1(111, 22)    <= sub_wire17(22);
	sub_wire1(111, 23)    <= sub_wire17(23);
	sub_wire1(111, 24)    <= sub_wire17(24);
	sub_wire1(111, 25)    <= sub_wire17(25);
	sub_wire1(111, 26)    <= sub_wire17(26);
	sub_wire1(111, 27)    <= sub_wire17(27);
	sub_wire1(111, 28)    <= sub_wire17(28);
	sub_wire1(111, 29)    <= sub_wire17(29);
	sub_wire1(111, 30)    <= sub_wire17(30);
	sub_wire1(111, 31)    <= sub_wire17(31);
	sub_wire1(110, 0)    <= sub_wire18(0);
	sub_wire1(110, 1)    <= sub_wire18(1);
	sub_wire1(110, 2)    <= sub_wire18(2);
	sub_wire1(110, 3)    <= sub_wire18(3);
	sub_wire1(110, 4)    <= sub_wire18(4);
	sub_wire1(110, 5)    <= sub_wire18(5);
	sub_wire1(110, 6)    <= sub_wire18(6);
	sub_wire1(110, 7)    <= sub_wire18(7);
	sub_wire1(110, 8)    <= sub_wire18(8);
	sub_wire1(110, 9)    <= sub_wire18(9);
	sub_wire1(110, 10)    <= sub_wire18(10);
	sub_wire1(110, 11)    <= sub_wire18(11);
	sub_wire1(110, 12)    <= sub_wire18(12);
	sub_wire1(110, 13)    <= sub_wire18(13);
	sub_wire1(110, 14)    <= sub_wire18(14);
	sub_wire1(110, 15)    <= sub_wire18(15);
	sub_wire1(110, 16)    <= sub_wire18(16);
	sub_wire1(110, 17)    <= sub_wire18(17);
	sub_wire1(110, 18)    <= sub_wire18(18);
	sub_wire1(110, 19)    <= sub_wire18(19);
	sub_wire1(110, 20)    <= sub_wire18(20);
	sub_wire1(110, 21)    <= sub_wire18(21);
	sub_wire1(110, 22)    <= sub_wire18(22);
	sub_wire1(110, 23)    <= sub_wire18(23);
	sub_wire1(110, 24)    <= sub_wire18(24);
	sub_wire1(110, 25)    <= sub_wire18(25);
	sub_wire1(110, 26)    <= sub_wire18(26);
	sub_wire1(110, 27)    <= sub_wire18(27);
	sub_wire1(110, 28)    <= sub_wire18(28);
	sub_wire1(110, 29)    <= sub_wire18(29);
	sub_wire1(110, 30)    <= sub_wire18(30);
	sub_wire1(110, 31)    <= sub_wire18(31);
	sub_wire1(109, 0)    <= sub_wire19(0);
	sub_wire1(109, 1)    <= sub_wire19(1);
	sub_wire1(109, 2)    <= sub_wire19(2);
	sub_wire1(109, 3)    <= sub_wire19(3);
	sub_wire1(109, 4)    <= sub_wire19(4);
	sub_wire1(109, 5)    <= sub_wire19(5);
	sub_wire1(109, 6)    <= sub_wire19(6);
	sub_wire1(109, 7)    <= sub_wire19(7);
	sub_wire1(109, 8)    <= sub_wire19(8);
	sub_wire1(109, 9)    <= sub_wire19(9);
	sub_wire1(109, 10)    <= sub_wire19(10);
	sub_wire1(109, 11)    <= sub_wire19(11);
	sub_wire1(109, 12)    <= sub_wire19(12);
	sub_wire1(109, 13)    <= sub_wire19(13);
	sub_wire1(109, 14)    <= sub_wire19(14);
	sub_wire1(109, 15)    <= sub_wire19(15);
	sub_wire1(109, 16)    <= sub_wire19(16);
	sub_wire1(109, 17)    <= sub_wire19(17);
	sub_wire1(109, 18)    <= sub_wire19(18);
	sub_wire1(109, 19)    <= sub_wire19(19);
	sub_wire1(109, 20)    <= sub_wire19(20);
	sub_wire1(109, 21)    <= sub_wire19(21);
	sub_wire1(109, 22)    <= sub_wire19(22);
	sub_wire1(109, 23)    <= sub_wire19(23);
	sub_wire1(109, 24)    <= sub_wire19(24);
	sub_wire1(109, 25)    <= sub_wire19(25);
	sub_wire1(109, 26)    <= sub_wire19(26);
	sub_wire1(109, 27)    <= sub_wire19(27);
	sub_wire1(109, 28)    <= sub_wire19(28);
	sub_wire1(109, 29)    <= sub_wire19(29);
	sub_wire1(109, 30)    <= sub_wire19(30);
	sub_wire1(109, 31)    <= sub_wire19(31);
	sub_wire1(108, 0)    <= sub_wire20(0);
	sub_wire1(108, 1)    <= sub_wire20(1);
	sub_wire1(108, 2)    <= sub_wire20(2);
	sub_wire1(108, 3)    <= sub_wire20(3);
	sub_wire1(108, 4)    <= sub_wire20(4);
	sub_wire1(108, 5)    <= sub_wire20(5);
	sub_wire1(108, 6)    <= sub_wire20(6);
	sub_wire1(108, 7)    <= sub_wire20(7);
	sub_wire1(108, 8)    <= sub_wire20(8);
	sub_wire1(108, 9)    <= sub_wire20(9);
	sub_wire1(108, 10)    <= sub_wire20(10);
	sub_wire1(108, 11)    <= sub_wire20(11);
	sub_wire1(108, 12)    <= sub_wire20(12);
	sub_wire1(108, 13)    <= sub_wire20(13);
	sub_wire1(108, 14)    <= sub_wire20(14);
	sub_wire1(108, 15)    <= sub_wire20(15);
	sub_wire1(108, 16)    <= sub_wire20(16);
	sub_wire1(108, 17)    <= sub_wire20(17);
	sub_wire1(108, 18)    <= sub_wire20(18);
	sub_wire1(108, 19)    <= sub_wire20(19);
	sub_wire1(108, 20)    <= sub_wire20(20);
	sub_wire1(108, 21)    <= sub_wire20(21);
	sub_wire1(108, 22)    <= sub_wire20(22);
	sub_wire1(108, 23)    <= sub_wire20(23);
	sub_wire1(108, 24)    <= sub_wire20(24);
	sub_wire1(108, 25)    <= sub_wire20(25);
	sub_wire1(108, 26)    <= sub_wire20(26);
	sub_wire1(108, 27)    <= sub_wire20(27);
	sub_wire1(108, 28)    <= sub_wire20(28);
	sub_wire1(108, 29)    <= sub_wire20(29);
	sub_wire1(108, 30)    <= sub_wire20(30);
	sub_wire1(108, 31)    <= sub_wire20(31);
	sub_wire1(107, 0)    <= sub_wire21(0);
	sub_wire1(107, 1)    <= sub_wire21(1);
	sub_wire1(107, 2)    <= sub_wire21(2);
	sub_wire1(107, 3)    <= sub_wire21(3);
	sub_wire1(107, 4)    <= sub_wire21(4);
	sub_wire1(107, 5)    <= sub_wire21(5);
	sub_wire1(107, 6)    <= sub_wire21(6);
	sub_wire1(107, 7)    <= sub_wire21(7);
	sub_wire1(107, 8)    <= sub_wire21(8);
	sub_wire1(107, 9)    <= sub_wire21(9);
	sub_wire1(107, 10)    <= sub_wire21(10);
	sub_wire1(107, 11)    <= sub_wire21(11);
	sub_wire1(107, 12)    <= sub_wire21(12);
	sub_wire1(107, 13)    <= sub_wire21(13);
	sub_wire1(107, 14)    <= sub_wire21(14);
	sub_wire1(107, 15)    <= sub_wire21(15);
	sub_wire1(107, 16)    <= sub_wire21(16);
	sub_wire1(107, 17)    <= sub_wire21(17);
	sub_wire1(107, 18)    <= sub_wire21(18);
	sub_wire1(107, 19)    <= sub_wire21(19);
	sub_wire1(107, 20)    <= sub_wire21(20);
	sub_wire1(107, 21)    <= sub_wire21(21);
	sub_wire1(107, 22)    <= sub_wire21(22);
	sub_wire1(107, 23)    <= sub_wire21(23);
	sub_wire1(107, 24)    <= sub_wire21(24);
	sub_wire1(107, 25)    <= sub_wire21(25);
	sub_wire1(107, 26)    <= sub_wire21(26);
	sub_wire1(107, 27)    <= sub_wire21(27);
	sub_wire1(107, 28)    <= sub_wire21(28);
	sub_wire1(107, 29)    <= sub_wire21(29);
	sub_wire1(107, 30)    <= sub_wire21(30);
	sub_wire1(107, 31)    <= sub_wire21(31);
	sub_wire1(106, 0)    <= sub_wire22(0);
	sub_wire1(106, 1)    <= sub_wire22(1);
	sub_wire1(106, 2)    <= sub_wire22(2);
	sub_wire1(106, 3)    <= sub_wire22(3);
	sub_wire1(106, 4)    <= sub_wire22(4);
	sub_wire1(106, 5)    <= sub_wire22(5);
	sub_wire1(106, 6)    <= sub_wire22(6);
	sub_wire1(106, 7)    <= sub_wire22(7);
	sub_wire1(106, 8)    <= sub_wire22(8);
	sub_wire1(106, 9)    <= sub_wire22(9);
	sub_wire1(106, 10)    <= sub_wire22(10);
	sub_wire1(106, 11)    <= sub_wire22(11);
	sub_wire1(106, 12)    <= sub_wire22(12);
	sub_wire1(106, 13)    <= sub_wire22(13);
	sub_wire1(106, 14)    <= sub_wire22(14);
	sub_wire1(106, 15)    <= sub_wire22(15);
	sub_wire1(106, 16)    <= sub_wire22(16);
	sub_wire1(106, 17)    <= sub_wire22(17);
	sub_wire1(106, 18)    <= sub_wire22(18);
	sub_wire1(106, 19)    <= sub_wire22(19);
	sub_wire1(106, 20)    <= sub_wire22(20);
	sub_wire1(106, 21)    <= sub_wire22(21);
	sub_wire1(106, 22)    <= sub_wire22(22);
	sub_wire1(106, 23)    <= sub_wire22(23);
	sub_wire1(106, 24)    <= sub_wire22(24);
	sub_wire1(106, 25)    <= sub_wire22(25);
	sub_wire1(106, 26)    <= sub_wire22(26);
	sub_wire1(106, 27)    <= sub_wire22(27);
	sub_wire1(106, 28)    <= sub_wire22(28);
	sub_wire1(106, 29)    <= sub_wire22(29);
	sub_wire1(106, 30)    <= sub_wire22(30);
	sub_wire1(106, 31)    <= sub_wire22(31);
	sub_wire1(105, 0)    <= sub_wire23(0);
	sub_wire1(105, 1)    <= sub_wire23(1);
	sub_wire1(105, 2)    <= sub_wire23(2);
	sub_wire1(105, 3)    <= sub_wire23(3);
	sub_wire1(105, 4)    <= sub_wire23(4);
	sub_wire1(105, 5)    <= sub_wire23(5);
	sub_wire1(105, 6)    <= sub_wire23(6);
	sub_wire1(105, 7)    <= sub_wire23(7);
	sub_wire1(105, 8)    <= sub_wire23(8);
	sub_wire1(105, 9)    <= sub_wire23(9);
	sub_wire1(105, 10)    <= sub_wire23(10);
	sub_wire1(105, 11)    <= sub_wire23(11);
	sub_wire1(105, 12)    <= sub_wire23(12);
	sub_wire1(105, 13)    <= sub_wire23(13);
	sub_wire1(105, 14)    <= sub_wire23(14);
	sub_wire1(105, 15)    <= sub_wire23(15);
	sub_wire1(105, 16)    <= sub_wire23(16);
	sub_wire1(105, 17)    <= sub_wire23(17);
	sub_wire1(105, 18)    <= sub_wire23(18);
	sub_wire1(105, 19)    <= sub_wire23(19);
	sub_wire1(105, 20)    <= sub_wire23(20);
	sub_wire1(105, 21)    <= sub_wire23(21);
	sub_wire1(105, 22)    <= sub_wire23(22);
	sub_wire1(105, 23)    <= sub_wire23(23);
	sub_wire1(105, 24)    <= sub_wire23(24);
	sub_wire1(105, 25)    <= sub_wire23(25);
	sub_wire1(105, 26)    <= sub_wire23(26);
	sub_wire1(105, 27)    <= sub_wire23(27);
	sub_wire1(105, 28)    <= sub_wire23(28);
	sub_wire1(105, 29)    <= sub_wire23(29);
	sub_wire1(105, 30)    <= sub_wire23(30);
	sub_wire1(105, 31)    <= sub_wire23(31);
	sub_wire1(104, 0)    <= sub_wire24(0);
	sub_wire1(104, 1)    <= sub_wire24(1);
	sub_wire1(104, 2)    <= sub_wire24(2);
	sub_wire1(104, 3)    <= sub_wire24(3);
	sub_wire1(104, 4)    <= sub_wire24(4);
	sub_wire1(104, 5)    <= sub_wire24(5);
	sub_wire1(104, 6)    <= sub_wire24(6);
	sub_wire1(104, 7)    <= sub_wire24(7);
	sub_wire1(104, 8)    <= sub_wire24(8);
	sub_wire1(104, 9)    <= sub_wire24(9);
	sub_wire1(104, 10)    <= sub_wire24(10);
	sub_wire1(104, 11)    <= sub_wire24(11);
	sub_wire1(104, 12)    <= sub_wire24(12);
	sub_wire1(104, 13)    <= sub_wire24(13);
	sub_wire1(104, 14)    <= sub_wire24(14);
	sub_wire1(104, 15)    <= sub_wire24(15);
	sub_wire1(104, 16)    <= sub_wire24(16);
	sub_wire1(104, 17)    <= sub_wire24(17);
	sub_wire1(104, 18)    <= sub_wire24(18);
	sub_wire1(104, 19)    <= sub_wire24(19);
	sub_wire1(104, 20)    <= sub_wire24(20);
	sub_wire1(104, 21)    <= sub_wire24(21);
	sub_wire1(104, 22)    <= sub_wire24(22);
	sub_wire1(104, 23)    <= sub_wire24(23);
	sub_wire1(104, 24)    <= sub_wire24(24);
	sub_wire1(104, 25)    <= sub_wire24(25);
	sub_wire1(104, 26)    <= sub_wire24(26);
	sub_wire1(104, 27)    <= sub_wire24(27);
	sub_wire1(104, 28)    <= sub_wire24(28);
	sub_wire1(104, 29)    <= sub_wire24(29);
	sub_wire1(104, 30)    <= sub_wire24(30);
	sub_wire1(104, 31)    <= sub_wire24(31);
	sub_wire1(103, 0)    <= sub_wire25(0);
	sub_wire1(103, 1)    <= sub_wire25(1);
	sub_wire1(103, 2)    <= sub_wire25(2);
	sub_wire1(103, 3)    <= sub_wire25(3);
	sub_wire1(103, 4)    <= sub_wire25(4);
	sub_wire1(103, 5)    <= sub_wire25(5);
	sub_wire1(103, 6)    <= sub_wire25(6);
	sub_wire1(103, 7)    <= sub_wire25(7);
	sub_wire1(103, 8)    <= sub_wire25(8);
	sub_wire1(103, 9)    <= sub_wire25(9);
	sub_wire1(103, 10)    <= sub_wire25(10);
	sub_wire1(103, 11)    <= sub_wire25(11);
	sub_wire1(103, 12)    <= sub_wire25(12);
	sub_wire1(103, 13)    <= sub_wire25(13);
	sub_wire1(103, 14)    <= sub_wire25(14);
	sub_wire1(103, 15)    <= sub_wire25(15);
	sub_wire1(103, 16)    <= sub_wire25(16);
	sub_wire1(103, 17)    <= sub_wire25(17);
	sub_wire1(103, 18)    <= sub_wire25(18);
	sub_wire1(103, 19)    <= sub_wire25(19);
	sub_wire1(103, 20)    <= sub_wire25(20);
	sub_wire1(103, 21)    <= sub_wire25(21);
	sub_wire1(103, 22)    <= sub_wire25(22);
	sub_wire1(103, 23)    <= sub_wire25(23);
	sub_wire1(103, 24)    <= sub_wire25(24);
	sub_wire1(103, 25)    <= sub_wire25(25);
	sub_wire1(103, 26)    <= sub_wire25(26);
	sub_wire1(103, 27)    <= sub_wire25(27);
	sub_wire1(103, 28)    <= sub_wire25(28);
	sub_wire1(103, 29)    <= sub_wire25(29);
	sub_wire1(103, 30)    <= sub_wire25(30);
	sub_wire1(103, 31)    <= sub_wire25(31);
	sub_wire1(102, 0)    <= sub_wire26(0);
	sub_wire1(102, 1)    <= sub_wire26(1);
	sub_wire1(102, 2)    <= sub_wire26(2);
	sub_wire1(102, 3)    <= sub_wire26(3);
	sub_wire1(102, 4)    <= sub_wire26(4);
	sub_wire1(102, 5)    <= sub_wire26(5);
	sub_wire1(102, 6)    <= sub_wire26(6);
	sub_wire1(102, 7)    <= sub_wire26(7);
	sub_wire1(102, 8)    <= sub_wire26(8);
	sub_wire1(102, 9)    <= sub_wire26(9);
	sub_wire1(102, 10)    <= sub_wire26(10);
	sub_wire1(102, 11)    <= sub_wire26(11);
	sub_wire1(102, 12)    <= sub_wire26(12);
	sub_wire1(102, 13)    <= sub_wire26(13);
	sub_wire1(102, 14)    <= sub_wire26(14);
	sub_wire1(102, 15)    <= sub_wire26(15);
	sub_wire1(102, 16)    <= sub_wire26(16);
	sub_wire1(102, 17)    <= sub_wire26(17);
	sub_wire1(102, 18)    <= sub_wire26(18);
	sub_wire1(102, 19)    <= sub_wire26(19);
	sub_wire1(102, 20)    <= sub_wire26(20);
	sub_wire1(102, 21)    <= sub_wire26(21);
	sub_wire1(102, 22)    <= sub_wire26(22);
	sub_wire1(102, 23)    <= sub_wire26(23);
	sub_wire1(102, 24)    <= sub_wire26(24);
	sub_wire1(102, 25)    <= sub_wire26(25);
	sub_wire1(102, 26)    <= sub_wire26(26);
	sub_wire1(102, 27)    <= sub_wire26(27);
	sub_wire1(102, 28)    <= sub_wire26(28);
	sub_wire1(102, 29)    <= sub_wire26(29);
	sub_wire1(102, 30)    <= sub_wire26(30);
	sub_wire1(102, 31)    <= sub_wire26(31);
	sub_wire1(101, 0)    <= sub_wire27(0);
	sub_wire1(101, 1)    <= sub_wire27(1);
	sub_wire1(101, 2)    <= sub_wire27(2);
	sub_wire1(101, 3)    <= sub_wire27(3);
	sub_wire1(101, 4)    <= sub_wire27(4);
	sub_wire1(101, 5)    <= sub_wire27(5);
	sub_wire1(101, 6)    <= sub_wire27(6);
	sub_wire1(101, 7)    <= sub_wire27(7);
	sub_wire1(101, 8)    <= sub_wire27(8);
	sub_wire1(101, 9)    <= sub_wire27(9);
	sub_wire1(101, 10)    <= sub_wire27(10);
	sub_wire1(101, 11)    <= sub_wire27(11);
	sub_wire1(101, 12)    <= sub_wire27(12);
	sub_wire1(101, 13)    <= sub_wire27(13);
	sub_wire1(101, 14)    <= sub_wire27(14);
	sub_wire1(101, 15)    <= sub_wire27(15);
	sub_wire1(101, 16)    <= sub_wire27(16);
	sub_wire1(101, 17)    <= sub_wire27(17);
	sub_wire1(101, 18)    <= sub_wire27(18);
	sub_wire1(101, 19)    <= sub_wire27(19);
	sub_wire1(101, 20)    <= sub_wire27(20);
	sub_wire1(101, 21)    <= sub_wire27(21);
	sub_wire1(101, 22)    <= sub_wire27(22);
	sub_wire1(101, 23)    <= sub_wire27(23);
	sub_wire1(101, 24)    <= sub_wire27(24);
	sub_wire1(101, 25)    <= sub_wire27(25);
	sub_wire1(101, 26)    <= sub_wire27(26);
	sub_wire1(101, 27)    <= sub_wire27(27);
	sub_wire1(101, 28)    <= sub_wire27(28);
	sub_wire1(101, 29)    <= sub_wire27(29);
	sub_wire1(101, 30)    <= sub_wire27(30);
	sub_wire1(101, 31)    <= sub_wire27(31);
	sub_wire1(100, 0)    <= sub_wire28(0);
	sub_wire1(100, 1)    <= sub_wire28(1);
	sub_wire1(100, 2)    <= sub_wire28(2);
	sub_wire1(100, 3)    <= sub_wire28(3);
	sub_wire1(100, 4)    <= sub_wire28(4);
	sub_wire1(100, 5)    <= sub_wire28(5);
	sub_wire1(100, 6)    <= sub_wire28(6);
	sub_wire1(100, 7)    <= sub_wire28(7);
	sub_wire1(100, 8)    <= sub_wire28(8);
	sub_wire1(100, 9)    <= sub_wire28(9);
	sub_wire1(100, 10)    <= sub_wire28(10);
	sub_wire1(100, 11)    <= sub_wire28(11);
	sub_wire1(100, 12)    <= sub_wire28(12);
	sub_wire1(100, 13)    <= sub_wire28(13);
	sub_wire1(100, 14)    <= sub_wire28(14);
	sub_wire1(100, 15)    <= sub_wire28(15);
	sub_wire1(100, 16)    <= sub_wire28(16);
	sub_wire1(100, 17)    <= sub_wire28(17);
	sub_wire1(100, 18)    <= sub_wire28(18);
	sub_wire1(100, 19)    <= sub_wire28(19);
	sub_wire1(100, 20)    <= sub_wire28(20);
	sub_wire1(100, 21)    <= sub_wire28(21);
	sub_wire1(100, 22)    <= sub_wire28(22);
	sub_wire1(100, 23)    <= sub_wire28(23);
	sub_wire1(100, 24)    <= sub_wire28(24);
	sub_wire1(100, 25)    <= sub_wire28(25);
	sub_wire1(100, 26)    <= sub_wire28(26);
	sub_wire1(100, 27)    <= sub_wire28(27);
	sub_wire1(100, 28)    <= sub_wire28(28);
	sub_wire1(100, 29)    <= sub_wire28(29);
	sub_wire1(100, 30)    <= sub_wire28(30);
	sub_wire1(100, 31)    <= sub_wire28(31);
	sub_wire1(99, 0)    <= sub_wire29(0);
	sub_wire1(99, 1)    <= sub_wire29(1);
	sub_wire1(99, 2)    <= sub_wire29(2);
	sub_wire1(99, 3)    <= sub_wire29(3);
	sub_wire1(99, 4)    <= sub_wire29(4);
	sub_wire1(99, 5)    <= sub_wire29(5);
	sub_wire1(99, 6)    <= sub_wire29(6);
	sub_wire1(99, 7)    <= sub_wire29(7);
	sub_wire1(99, 8)    <= sub_wire29(8);
	sub_wire1(99, 9)    <= sub_wire29(9);
	sub_wire1(99, 10)    <= sub_wire29(10);
	sub_wire1(99, 11)    <= sub_wire29(11);
	sub_wire1(99, 12)    <= sub_wire29(12);
	sub_wire1(99, 13)    <= sub_wire29(13);
	sub_wire1(99, 14)    <= sub_wire29(14);
	sub_wire1(99, 15)    <= sub_wire29(15);
	sub_wire1(99, 16)    <= sub_wire29(16);
	sub_wire1(99, 17)    <= sub_wire29(17);
	sub_wire1(99, 18)    <= sub_wire29(18);
	sub_wire1(99, 19)    <= sub_wire29(19);
	sub_wire1(99, 20)    <= sub_wire29(20);
	sub_wire1(99, 21)    <= sub_wire29(21);
	sub_wire1(99, 22)    <= sub_wire29(22);
	sub_wire1(99, 23)    <= sub_wire29(23);
	sub_wire1(99, 24)    <= sub_wire29(24);
	sub_wire1(99, 25)    <= sub_wire29(25);
	sub_wire1(99, 26)    <= sub_wire29(26);
	sub_wire1(99, 27)    <= sub_wire29(27);
	sub_wire1(99, 28)    <= sub_wire29(28);
	sub_wire1(99, 29)    <= sub_wire29(29);
	sub_wire1(99, 30)    <= sub_wire29(30);
	sub_wire1(99, 31)    <= sub_wire29(31);
	sub_wire1(98, 0)    <= sub_wire30(0);
	sub_wire1(98, 1)    <= sub_wire30(1);
	sub_wire1(98, 2)    <= sub_wire30(2);
	sub_wire1(98, 3)    <= sub_wire30(3);
	sub_wire1(98, 4)    <= sub_wire30(4);
	sub_wire1(98, 5)    <= sub_wire30(5);
	sub_wire1(98, 6)    <= sub_wire30(6);
	sub_wire1(98, 7)    <= sub_wire30(7);
	sub_wire1(98, 8)    <= sub_wire30(8);
	sub_wire1(98, 9)    <= sub_wire30(9);
	sub_wire1(98, 10)    <= sub_wire30(10);
	sub_wire1(98, 11)    <= sub_wire30(11);
	sub_wire1(98, 12)    <= sub_wire30(12);
	sub_wire1(98, 13)    <= sub_wire30(13);
	sub_wire1(98, 14)    <= sub_wire30(14);
	sub_wire1(98, 15)    <= sub_wire30(15);
	sub_wire1(98, 16)    <= sub_wire30(16);
	sub_wire1(98, 17)    <= sub_wire30(17);
	sub_wire1(98, 18)    <= sub_wire30(18);
	sub_wire1(98, 19)    <= sub_wire30(19);
	sub_wire1(98, 20)    <= sub_wire30(20);
	sub_wire1(98, 21)    <= sub_wire30(21);
	sub_wire1(98, 22)    <= sub_wire30(22);
	sub_wire1(98, 23)    <= sub_wire30(23);
	sub_wire1(98, 24)    <= sub_wire30(24);
	sub_wire1(98, 25)    <= sub_wire30(25);
	sub_wire1(98, 26)    <= sub_wire30(26);
	sub_wire1(98, 27)    <= sub_wire30(27);
	sub_wire1(98, 28)    <= sub_wire30(28);
	sub_wire1(98, 29)    <= sub_wire30(29);
	sub_wire1(98, 30)    <= sub_wire30(30);
	sub_wire1(98, 31)    <= sub_wire30(31);
	sub_wire1(97, 0)    <= sub_wire31(0);
	sub_wire1(97, 1)    <= sub_wire31(1);
	sub_wire1(97, 2)    <= sub_wire31(2);
	sub_wire1(97, 3)    <= sub_wire31(3);
	sub_wire1(97, 4)    <= sub_wire31(4);
	sub_wire1(97, 5)    <= sub_wire31(5);
	sub_wire1(97, 6)    <= sub_wire31(6);
	sub_wire1(97, 7)    <= sub_wire31(7);
	sub_wire1(97, 8)    <= sub_wire31(8);
	sub_wire1(97, 9)    <= sub_wire31(9);
	sub_wire1(97, 10)    <= sub_wire31(10);
	sub_wire1(97, 11)    <= sub_wire31(11);
	sub_wire1(97, 12)    <= sub_wire31(12);
	sub_wire1(97, 13)    <= sub_wire31(13);
	sub_wire1(97, 14)    <= sub_wire31(14);
	sub_wire1(97, 15)    <= sub_wire31(15);
	sub_wire1(97, 16)    <= sub_wire31(16);
	sub_wire1(97, 17)    <= sub_wire31(17);
	sub_wire1(97, 18)    <= sub_wire31(18);
	sub_wire1(97, 19)    <= sub_wire31(19);
	sub_wire1(97, 20)    <= sub_wire31(20);
	sub_wire1(97, 21)    <= sub_wire31(21);
	sub_wire1(97, 22)    <= sub_wire31(22);
	sub_wire1(97, 23)    <= sub_wire31(23);
	sub_wire1(97, 24)    <= sub_wire31(24);
	sub_wire1(97, 25)    <= sub_wire31(25);
	sub_wire1(97, 26)    <= sub_wire31(26);
	sub_wire1(97, 27)    <= sub_wire31(27);
	sub_wire1(97, 28)    <= sub_wire31(28);
	sub_wire1(97, 29)    <= sub_wire31(29);
	sub_wire1(97, 30)    <= sub_wire31(30);
	sub_wire1(97, 31)    <= sub_wire31(31);
	sub_wire1(96, 0)    <= sub_wire32(0);
	sub_wire1(96, 1)    <= sub_wire32(1);
	sub_wire1(96, 2)    <= sub_wire32(2);
	sub_wire1(96, 3)    <= sub_wire32(3);
	sub_wire1(96, 4)    <= sub_wire32(4);
	sub_wire1(96, 5)    <= sub_wire32(5);
	sub_wire1(96, 6)    <= sub_wire32(6);
	sub_wire1(96, 7)    <= sub_wire32(7);
	sub_wire1(96, 8)    <= sub_wire32(8);
	sub_wire1(96, 9)    <= sub_wire32(9);
	sub_wire1(96, 10)    <= sub_wire32(10);
	sub_wire1(96, 11)    <= sub_wire32(11);
	sub_wire1(96, 12)    <= sub_wire32(12);
	sub_wire1(96, 13)    <= sub_wire32(13);
	sub_wire1(96, 14)    <= sub_wire32(14);
	sub_wire1(96, 15)    <= sub_wire32(15);
	sub_wire1(96, 16)    <= sub_wire32(16);
	sub_wire1(96, 17)    <= sub_wire32(17);
	sub_wire1(96, 18)    <= sub_wire32(18);
	sub_wire1(96, 19)    <= sub_wire32(19);
	sub_wire1(96, 20)    <= sub_wire32(20);
	sub_wire1(96, 21)    <= sub_wire32(21);
	sub_wire1(96, 22)    <= sub_wire32(22);
	sub_wire1(96, 23)    <= sub_wire32(23);
	sub_wire1(96, 24)    <= sub_wire32(24);
	sub_wire1(96, 25)    <= sub_wire32(25);
	sub_wire1(96, 26)    <= sub_wire32(26);
	sub_wire1(96, 27)    <= sub_wire32(27);
	sub_wire1(96, 28)    <= sub_wire32(28);
	sub_wire1(96, 29)    <= sub_wire32(29);
	sub_wire1(96, 30)    <= sub_wire32(30);
	sub_wire1(96, 31)    <= sub_wire32(31);
	sub_wire1(95, 0)    <= sub_wire33(0);
	sub_wire1(95, 1)    <= sub_wire33(1);
	sub_wire1(95, 2)    <= sub_wire33(2);
	sub_wire1(95, 3)    <= sub_wire33(3);
	sub_wire1(95, 4)    <= sub_wire33(4);
	sub_wire1(95, 5)    <= sub_wire33(5);
	sub_wire1(95, 6)    <= sub_wire33(6);
	sub_wire1(95, 7)    <= sub_wire33(7);
	sub_wire1(95, 8)    <= sub_wire33(8);
	sub_wire1(95, 9)    <= sub_wire33(9);
	sub_wire1(95, 10)    <= sub_wire33(10);
	sub_wire1(95, 11)    <= sub_wire33(11);
	sub_wire1(95, 12)    <= sub_wire33(12);
	sub_wire1(95, 13)    <= sub_wire33(13);
	sub_wire1(95, 14)    <= sub_wire33(14);
	sub_wire1(95, 15)    <= sub_wire33(15);
	sub_wire1(95, 16)    <= sub_wire33(16);
	sub_wire1(95, 17)    <= sub_wire33(17);
	sub_wire1(95, 18)    <= sub_wire33(18);
	sub_wire1(95, 19)    <= sub_wire33(19);
	sub_wire1(95, 20)    <= sub_wire33(20);
	sub_wire1(95, 21)    <= sub_wire33(21);
	sub_wire1(95, 22)    <= sub_wire33(22);
	sub_wire1(95, 23)    <= sub_wire33(23);
	sub_wire1(95, 24)    <= sub_wire33(24);
	sub_wire1(95, 25)    <= sub_wire33(25);
	sub_wire1(95, 26)    <= sub_wire33(26);
	sub_wire1(95, 27)    <= sub_wire33(27);
	sub_wire1(95, 28)    <= sub_wire33(28);
	sub_wire1(95, 29)    <= sub_wire33(29);
	sub_wire1(95, 30)    <= sub_wire33(30);
	sub_wire1(95, 31)    <= sub_wire33(31);
	sub_wire1(94, 0)    <= sub_wire34(0);
	sub_wire1(94, 1)    <= sub_wire34(1);
	sub_wire1(94, 2)    <= sub_wire34(2);
	sub_wire1(94, 3)    <= sub_wire34(3);
	sub_wire1(94, 4)    <= sub_wire34(4);
	sub_wire1(94, 5)    <= sub_wire34(5);
	sub_wire1(94, 6)    <= sub_wire34(6);
	sub_wire1(94, 7)    <= sub_wire34(7);
	sub_wire1(94, 8)    <= sub_wire34(8);
	sub_wire1(94, 9)    <= sub_wire34(9);
	sub_wire1(94, 10)    <= sub_wire34(10);
	sub_wire1(94, 11)    <= sub_wire34(11);
	sub_wire1(94, 12)    <= sub_wire34(12);
	sub_wire1(94, 13)    <= sub_wire34(13);
	sub_wire1(94, 14)    <= sub_wire34(14);
	sub_wire1(94, 15)    <= sub_wire34(15);
	sub_wire1(94, 16)    <= sub_wire34(16);
	sub_wire1(94, 17)    <= sub_wire34(17);
	sub_wire1(94, 18)    <= sub_wire34(18);
	sub_wire1(94, 19)    <= sub_wire34(19);
	sub_wire1(94, 20)    <= sub_wire34(20);
	sub_wire1(94, 21)    <= sub_wire34(21);
	sub_wire1(94, 22)    <= sub_wire34(22);
	sub_wire1(94, 23)    <= sub_wire34(23);
	sub_wire1(94, 24)    <= sub_wire34(24);
	sub_wire1(94, 25)    <= sub_wire34(25);
	sub_wire1(94, 26)    <= sub_wire34(26);
	sub_wire1(94, 27)    <= sub_wire34(27);
	sub_wire1(94, 28)    <= sub_wire34(28);
	sub_wire1(94, 29)    <= sub_wire34(29);
	sub_wire1(94, 30)    <= sub_wire34(30);
	sub_wire1(94, 31)    <= sub_wire34(31);
	sub_wire1(93, 0)    <= sub_wire35(0);
	sub_wire1(93, 1)    <= sub_wire35(1);
	sub_wire1(93, 2)    <= sub_wire35(2);
	sub_wire1(93, 3)    <= sub_wire35(3);
	sub_wire1(93, 4)    <= sub_wire35(4);
	sub_wire1(93, 5)    <= sub_wire35(5);
	sub_wire1(93, 6)    <= sub_wire35(6);
	sub_wire1(93, 7)    <= sub_wire35(7);
	sub_wire1(93, 8)    <= sub_wire35(8);
	sub_wire1(93, 9)    <= sub_wire35(9);
	sub_wire1(93, 10)    <= sub_wire35(10);
	sub_wire1(93, 11)    <= sub_wire35(11);
	sub_wire1(93, 12)    <= sub_wire35(12);
	sub_wire1(93, 13)    <= sub_wire35(13);
	sub_wire1(93, 14)    <= sub_wire35(14);
	sub_wire1(93, 15)    <= sub_wire35(15);
	sub_wire1(93, 16)    <= sub_wire35(16);
	sub_wire1(93, 17)    <= sub_wire35(17);
	sub_wire1(93, 18)    <= sub_wire35(18);
	sub_wire1(93, 19)    <= sub_wire35(19);
	sub_wire1(93, 20)    <= sub_wire35(20);
	sub_wire1(93, 21)    <= sub_wire35(21);
	sub_wire1(93, 22)    <= sub_wire35(22);
	sub_wire1(93, 23)    <= sub_wire35(23);
	sub_wire1(93, 24)    <= sub_wire35(24);
	sub_wire1(93, 25)    <= sub_wire35(25);
	sub_wire1(93, 26)    <= sub_wire35(26);
	sub_wire1(93, 27)    <= sub_wire35(27);
	sub_wire1(93, 28)    <= sub_wire35(28);
	sub_wire1(93, 29)    <= sub_wire35(29);
	sub_wire1(93, 30)    <= sub_wire35(30);
	sub_wire1(93, 31)    <= sub_wire35(31);
	sub_wire1(92, 0)    <= sub_wire36(0);
	sub_wire1(92, 1)    <= sub_wire36(1);
	sub_wire1(92, 2)    <= sub_wire36(2);
	sub_wire1(92, 3)    <= sub_wire36(3);
	sub_wire1(92, 4)    <= sub_wire36(4);
	sub_wire1(92, 5)    <= sub_wire36(5);
	sub_wire1(92, 6)    <= sub_wire36(6);
	sub_wire1(92, 7)    <= sub_wire36(7);
	sub_wire1(92, 8)    <= sub_wire36(8);
	sub_wire1(92, 9)    <= sub_wire36(9);
	sub_wire1(92, 10)    <= sub_wire36(10);
	sub_wire1(92, 11)    <= sub_wire36(11);
	sub_wire1(92, 12)    <= sub_wire36(12);
	sub_wire1(92, 13)    <= sub_wire36(13);
	sub_wire1(92, 14)    <= sub_wire36(14);
	sub_wire1(92, 15)    <= sub_wire36(15);
	sub_wire1(92, 16)    <= sub_wire36(16);
	sub_wire1(92, 17)    <= sub_wire36(17);
	sub_wire1(92, 18)    <= sub_wire36(18);
	sub_wire1(92, 19)    <= sub_wire36(19);
	sub_wire1(92, 20)    <= sub_wire36(20);
	sub_wire1(92, 21)    <= sub_wire36(21);
	sub_wire1(92, 22)    <= sub_wire36(22);
	sub_wire1(92, 23)    <= sub_wire36(23);
	sub_wire1(92, 24)    <= sub_wire36(24);
	sub_wire1(92, 25)    <= sub_wire36(25);
	sub_wire1(92, 26)    <= sub_wire36(26);
	sub_wire1(92, 27)    <= sub_wire36(27);
	sub_wire1(92, 28)    <= sub_wire36(28);
	sub_wire1(92, 29)    <= sub_wire36(29);
	sub_wire1(92, 30)    <= sub_wire36(30);
	sub_wire1(92, 31)    <= sub_wire36(31);
	sub_wire1(91, 0)    <= sub_wire37(0);
	sub_wire1(91, 1)    <= sub_wire37(1);
	sub_wire1(91, 2)    <= sub_wire37(2);
	sub_wire1(91, 3)    <= sub_wire37(3);
	sub_wire1(91, 4)    <= sub_wire37(4);
	sub_wire1(91, 5)    <= sub_wire37(5);
	sub_wire1(91, 6)    <= sub_wire37(6);
	sub_wire1(91, 7)    <= sub_wire37(7);
	sub_wire1(91, 8)    <= sub_wire37(8);
	sub_wire1(91, 9)    <= sub_wire37(9);
	sub_wire1(91, 10)    <= sub_wire37(10);
	sub_wire1(91, 11)    <= sub_wire37(11);
	sub_wire1(91, 12)    <= sub_wire37(12);
	sub_wire1(91, 13)    <= sub_wire37(13);
	sub_wire1(91, 14)    <= sub_wire37(14);
	sub_wire1(91, 15)    <= sub_wire37(15);
	sub_wire1(91, 16)    <= sub_wire37(16);
	sub_wire1(91, 17)    <= sub_wire37(17);
	sub_wire1(91, 18)    <= sub_wire37(18);
	sub_wire1(91, 19)    <= sub_wire37(19);
	sub_wire1(91, 20)    <= sub_wire37(20);
	sub_wire1(91, 21)    <= sub_wire37(21);
	sub_wire1(91, 22)    <= sub_wire37(22);
	sub_wire1(91, 23)    <= sub_wire37(23);
	sub_wire1(91, 24)    <= sub_wire37(24);
	sub_wire1(91, 25)    <= sub_wire37(25);
	sub_wire1(91, 26)    <= sub_wire37(26);
	sub_wire1(91, 27)    <= sub_wire37(27);
	sub_wire1(91, 28)    <= sub_wire37(28);
	sub_wire1(91, 29)    <= sub_wire37(29);
	sub_wire1(91, 30)    <= sub_wire37(30);
	sub_wire1(91, 31)    <= sub_wire37(31);
	sub_wire1(90, 0)    <= sub_wire38(0);
	sub_wire1(90, 1)    <= sub_wire38(1);
	sub_wire1(90, 2)    <= sub_wire38(2);
	sub_wire1(90, 3)    <= sub_wire38(3);
	sub_wire1(90, 4)    <= sub_wire38(4);
	sub_wire1(90, 5)    <= sub_wire38(5);
	sub_wire1(90, 6)    <= sub_wire38(6);
	sub_wire1(90, 7)    <= sub_wire38(7);
	sub_wire1(90, 8)    <= sub_wire38(8);
	sub_wire1(90, 9)    <= sub_wire38(9);
	sub_wire1(90, 10)    <= sub_wire38(10);
	sub_wire1(90, 11)    <= sub_wire38(11);
	sub_wire1(90, 12)    <= sub_wire38(12);
	sub_wire1(90, 13)    <= sub_wire38(13);
	sub_wire1(90, 14)    <= sub_wire38(14);
	sub_wire1(90, 15)    <= sub_wire38(15);
	sub_wire1(90, 16)    <= sub_wire38(16);
	sub_wire1(90, 17)    <= sub_wire38(17);
	sub_wire1(90, 18)    <= sub_wire38(18);
	sub_wire1(90, 19)    <= sub_wire38(19);
	sub_wire1(90, 20)    <= sub_wire38(20);
	sub_wire1(90, 21)    <= sub_wire38(21);
	sub_wire1(90, 22)    <= sub_wire38(22);
	sub_wire1(90, 23)    <= sub_wire38(23);
	sub_wire1(90, 24)    <= sub_wire38(24);
	sub_wire1(90, 25)    <= sub_wire38(25);
	sub_wire1(90, 26)    <= sub_wire38(26);
	sub_wire1(90, 27)    <= sub_wire38(27);
	sub_wire1(90, 28)    <= sub_wire38(28);
	sub_wire1(90, 29)    <= sub_wire38(29);
	sub_wire1(90, 30)    <= sub_wire38(30);
	sub_wire1(90, 31)    <= sub_wire38(31);
	sub_wire1(89, 0)    <= sub_wire39(0);
	sub_wire1(89, 1)    <= sub_wire39(1);
	sub_wire1(89, 2)    <= sub_wire39(2);
	sub_wire1(89, 3)    <= sub_wire39(3);
	sub_wire1(89, 4)    <= sub_wire39(4);
	sub_wire1(89, 5)    <= sub_wire39(5);
	sub_wire1(89, 6)    <= sub_wire39(6);
	sub_wire1(89, 7)    <= sub_wire39(7);
	sub_wire1(89, 8)    <= sub_wire39(8);
	sub_wire1(89, 9)    <= sub_wire39(9);
	sub_wire1(89, 10)    <= sub_wire39(10);
	sub_wire1(89, 11)    <= sub_wire39(11);
	sub_wire1(89, 12)    <= sub_wire39(12);
	sub_wire1(89, 13)    <= sub_wire39(13);
	sub_wire1(89, 14)    <= sub_wire39(14);
	sub_wire1(89, 15)    <= sub_wire39(15);
	sub_wire1(89, 16)    <= sub_wire39(16);
	sub_wire1(89, 17)    <= sub_wire39(17);
	sub_wire1(89, 18)    <= sub_wire39(18);
	sub_wire1(89, 19)    <= sub_wire39(19);
	sub_wire1(89, 20)    <= sub_wire39(20);
	sub_wire1(89, 21)    <= sub_wire39(21);
	sub_wire1(89, 22)    <= sub_wire39(22);
	sub_wire1(89, 23)    <= sub_wire39(23);
	sub_wire1(89, 24)    <= sub_wire39(24);
	sub_wire1(89, 25)    <= sub_wire39(25);
	sub_wire1(89, 26)    <= sub_wire39(26);
	sub_wire1(89, 27)    <= sub_wire39(27);
	sub_wire1(89, 28)    <= sub_wire39(28);
	sub_wire1(89, 29)    <= sub_wire39(29);
	sub_wire1(89, 30)    <= sub_wire39(30);
	sub_wire1(89, 31)    <= sub_wire39(31);
	sub_wire1(88, 0)    <= sub_wire40(0);
	sub_wire1(88, 1)    <= sub_wire40(1);
	sub_wire1(88, 2)    <= sub_wire40(2);
	sub_wire1(88, 3)    <= sub_wire40(3);
	sub_wire1(88, 4)    <= sub_wire40(4);
	sub_wire1(88, 5)    <= sub_wire40(5);
	sub_wire1(88, 6)    <= sub_wire40(6);
	sub_wire1(88, 7)    <= sub_wire40(7);
	sub_wire1(88, 8)    <= sub_wire40(8);
	sub_wire1(88, 9)    <= sub_wire40(9);
	sub_wire1(88, 10)    <= sub_wire40(10);
	sub_wire1(88, 11)    <= sub_wire40(11);
	sub_wire1(88, 12)    <= sub_wire40(12);
	sub_wire1(88, 13)    <= sub_wire40(13);
	sub_wire1(88, 14)    <= sub_wire40(14);
	sub_wire1(88, 15)    <= sub_wire40(15);
	sub_wire1(88, 16)    <= sub_wire40(16);
	sub_wire1(88, 17)    <= sub_wire40(17);
	sub_wire1(88, 18)    <= sub_wire40(18);
	sub_wire1(88, 19)    <= sub_wire40(19);
	sub_wire1(88, 20)    <= sub_wire40(20);
	sub_wire1(88, 21)    <= sub_wire40(21);
	sub_wire1(88, 22)    <= sub_wire40(22);
	sub_wire1(88, 23)    <= sub_wire40(23);
	sub_wire1(88, 24)    <= sub_wire40(24);
	sub_wire1(88, 25)    <= sub_wire40(25);
	sub_wire1(88, 26)    <= sub_wire40(26);
	sub_wire1(88, 27)    <= sub_wire40(27);
	sub_wire1(88, 28)    <= sub_wire40(28);
	sub_wire1(88, 29)    <= sub_wire40(29);
	sub_wire1(88, 30)    <= sub_wire40(30);
	sub_wire1(88, 31)    <= sub_wire40(31);
	sub_wire1(87, 0)    <= sub_wire41(0);
	sub_wire1(87, 1)    <= sub_wire41(1);
	sub_wire1(87, 2)    <= sub_wire41(2);
	sub_wire1(87, 3)    <= sub_wire41(3);
	sub_wire1(87, 4)    <= sub_wire41(4);
	sub_wire1(87, 5)    <= sub_wire41(5);
	sub_wire1(87, 6)    <= sub_wire41(6);
	sub_wire1(87, 7)    <= sub_wire41(7);
	sub_wire1(87, 8)    <= sub_wire41(8);
	sub_wire1(87, 9)    <= sub_wire41(9);
	sub_wire1(87, 10)    <= sub_wire41(10);
	sub_wire1(87, 11)    <= sub_wire41(11);
	sub_wire1(87, 12)    <= sub_wire41(12);
	sub_wire1(87, 13)    <= sub_wire41(13);
	sub_wire1(87, 14)    <= sub_wire41(14);
	sub_wire1(87, 15)    <= sub_wire41(15);
	sub_wire1(87, 16)    <= sub_wire41(16);
	sub_wire1(87, 17)    <= sub_wire41(17);
	sub_wire1(87, 18)    <= sub_wire41(18);
	sub_wire1(87, 19)    <= sub_wire41(19);
	sub_wire1(87, 20)    <= sub_wire41(20);
	sub_wire1(87, 21)    <= sub_wire41(21);
	sub_wire1(87, 22)    <= sub_wire41(22);
	sub_wire1(87, 23)    <= sub_wire41(23);
	sub_wire1(87, 24)    <= sub_wire41(24);
	sub_wire1(87, 25)    <= sub_wire41(25);
	sub_wire1(87, 26)    <= sub_wire41(26);
	sub_wire1(87, 27)    <= sub_wire41(27);
	sub_wire1(87, 28)    <= sub_wire41(28);
	sub_wire1(87, 29)    <= sub_wire41(29);
	sub_wire1(87, 30)    <= sub_wire41(30);
	sub_wire1(87, 31)    <= sub_wire41(31);
	sub_wire1(86, 0)    <= sub_wire42(0);
	sub_wire1(86, 1)    <= sub_wire42(1);
	sub_wire1(86, 2)    <= sub_wire42(2);
	sub_wire1(86, 3)    <= sub_wire42(3);
	sub_wire1(86, 4)    <= sub_wire42(4);
	sub_wire1(86, 5)    <= sub_wire42(5);
	sub_wire1(86, 6)    <= sub_wire42(6);
	sub_wire1(86, 7)    <= sub_wire42(7);
	sub_wire1(86, 8)    <= sub_wire42(8);
	sub_wire1(86, 9)    <= sub_wire42(9);
	sub_wire1(86, 10)    <= sub_wire42(10);
	sub_wire1(86, 11)    <= sub_wire42(11);
	sub_wire1(86, 12)    <= sub_wire42(12);
	sub_wire1(86, 13)    <= sub_wire42(13);
	sub_wire1(86, 14)    <= sub_wire42(14);
	sub_wire1(86, 15)    <= sub_wire42(15);
	sub_wire1(86, 16)    <= sub_wire42(16);
	sub_wire1(86, 17)    <= sub_wire42(17);
	sub_wire1(86, 18)    <= sub_wire42(18);
	sub_wire1(86, 19)    <= sub_wire42(19);
	sub_wire1(86, 20)    <= sub_wire42(20);
	sub_wire1(86, 21)    <= sub_wire42(21);
	sub_wire1(86, 22)    <= sub_wire42(22);
	sub_wire1(86, 23)    <= sub_wire42(23);
	sub_wire1(86, 24)    <= sub_wire42(24);
	sub_wire1(86, 25)    <= sub_wire42(25);
	sub_wire1(86, 26)    <= sub_wire42(26);
	sub_wire1(86, 27)    <= sub_wire42(27);
	sub_wire1(86, 28)    <= sub_wire42(28);
	sub_wire1(86, 29)    <= sub_wire42(29);
	sub_wire1(86, 30)    <= sub_wire42(30);
	sub_wire1(86, 31)    <= sub_wire42(31);
	sub_wire1(85, 0)    <= sub_wire43(0);
	sub_wire1(85, 1)    <= sub_wire43(1);
	sub_wire1(85, 2)    <= sub_wire43(2);
	sub_wire1(85, 3)    <= sub_wire43(3);
	sub_wire1(85, 4)    <= sub_wire43(4);
	sub_wire1(85, 5)    <= sub_wire43(5);
	sub_wire1(85, 6)    <= sub_wire43(6);
	sub_wire1(85, 7)    <= sub_wire43(7);
	sub_wire1(85, 8)    <= sub_wire43(8);
	sub_wire1(85, 9)    <= sub_wire43(9);
	sub_wire1(85, 10)    <= sub_wire43(10);
	sub_wire1(85, 11)    <= sub_wire43(11);
	sub_wire1(85, 12)    <= sub_wire43(12);
	sub_wire1(85, 13)    <= sub_wire43(13);
	sub_wire1(85, 14)    <= sub_wire43(14);
	sub_wire1(85, 15)    <= sub_wire43(15);
	sub_wire1(85, 16)    <= sub_wire43(16);
	sub_wire1(85, 17)    <= sub_wire43(17);
	sub_wire1(85, 18)    <= sub_wire43(18);
	sub_wire1(85, 19)    <= sub_wire43(19);
	sub_wire1(85, 20)    <= sub_wire43(20);
	sub_wire1(85, 21)    <= sub_wire43(21);
	sub_wire1(85, 22)    <= sub_wire43(22);
	sub_wire1(85, 23)    <= sub_wire43(23);
	sub_wire1(85, 24)    <= sub_wire43(24);
	sub_wire1(85, 25)    <= sub_wire43(25);
	sub_wire1(85, 26)    <= sub_wire43(26);
	sub_wire1(85, 27)    <= sub_wire43(27);
	sub_wire1(85, 28)    <= sub_wire43(28);
	sub_wire1(85, 29)    <= sub_wire43(29);
	sub_wire1(85, 30)    <= sub_wire43(30);
	sub_wire1(85, 31)    <= sub_wire43(31);
	sub_wire1(84, 0)    <= sub_wire44(0);
	sub_wire1(84, 1)    <= sub_wire44(1);
	sub_wire1(84, 2)    <= sub_wire44(2);
	sub_wire1(84, 3)    <= sub_wire44(3);
	sub_wire1(84, 4)    <= sub_wire44(4);
	sub_wire1(84, 5)    <= sub_wire44(5);
	sub_wire1(84, 6)    <= sub_wire44(6);
	sub_wire1(84, 7)    <= sub_wire44(7);
	sub_wire1(84, 8)    <= sub_wire44(8);
	sub_wire1(84, 9)    <= sub_wire44(9);
	sub_wire1(84, 10)    <= sub_wire44(10);
	sub_wire1(84, 11)    <= sub_wire44(11);
	sub_wire1(84, 12)    <= sub_wire44(12);
	sub_wire1(84, 13)    <= sub_wire44(13);
	sub_wire1(84, 14)    <= sub_wire44(14);
	sub_wire1(84, 15)    <= sub_wire44(15);
	sub_wire1(84, 16)    <= sub_wire44(16);
	sub_wire1(84, 17)    <= sub_wire44(17);
	sub_wire1(84, 18)    <= sub_wire44(18);
	sub_wire1(84, 19)    <= sub_wire44(19);
	sub_wire1(84, 20)    <= sub_wire44(20);
	sub_wire1(84, 21)    <= sub_wire44(21);
	sub_wire1(84, 22)    <= sub_wire44(22);
	sub_wire1(84, 23)    <= sub_wire44(23);
	sub_wire1(84, 24)    <= sub_wire44(24);
	sub_wire1(84, 25)    <= sub_wire44(25);
	sub_wire1(84, 26)    <= sub_wire44(26);
	sub_wire1(84, 27)    <= sub_wire44(27);
	sub_wire1(84, 28)    <= sub_wire44(28);
	sub_wire1(84, 29)    <= sub_wire44(29);
	sub_wire1(84, 30)    <= sub_wire44(30);
	sub_wire1(84, 31)    <= sub_wire44(31);
	sub_wire1(83, 0)    <= sub_wire45(0);
	sub_wire1(83, 1)    <= sub_wire45(1);
	sub_wire1(83, 2)    <= sub_wire45(2);
	sub_wire1(83, 3)    <= sub_wire45(3);
	sub_wire1(83, 4)    <= sub_wire45(4);
	sub_wire1(83, 5)    <= sub_wire45(5);
	sub_wire1(83, 6)    <= sub_wire45(6);
	sub_wire1(83, 7)    <= sub_wire45(7);
	sub_wire1(83, 8)    <= sub_wire45(8);
	sub_wire1(83, 9)    <= sub_wire45(9);
	sub_wire1(83, 10)    <= sub_wire45(10);
	sub_wire1(83, 11)    <= sub_wire45(11);
	sub_wire1(83, 12)    <= sub_wire45(12);
	sub_wire1(83, 13)    <= sub_wire45(13);
	sub_wire1(83, 14)    <= sub_wire45(14);
	sub_wire1(83, 15)    <= sub_wire45(15);
	sub_wire1(83, 16)    <= sub_wire45(16);
	sub_wire1(83, 17)    <= sub_wire45(17);
	sub_wire1(83, 18)    <= sub_wire45(18);
	sub_wire1(83, 19)    <= sub_wire45(19);
	sub_wire1(83, 20)    <= sub_wire45(20);
	sub_wire1(83, 21)    <= sub_wire45(21);
	sub_wire1(83, 22)    <= sub_wire45(22);
	sub_wire1(83, 23)    <= sub_wire45(23);
	sub_wire1(83, 24)    <= sub_wire45(24);
	sub_wire1(83, 25)    <= sub_wire45(25);
	sub_wire1(83, 26)    <= sub_wire45(26);
	sub_wire1(83, 27)    <= sub_wire45(27);
	sub_wire1(83, 28)    <= sub_wire45(28);
	sub_wire1(83, 29)    <= sub_wire45(29);
	sub_wire1(83, 30)    <= sub_wire45(30);
	sub_wire1(83, 31)    <= sub_wire45(31);
	sub_wire1(82, 0)    <= sub_wire46(0);
	sub_wire1(82, 1)    <= sub_wire46(1);
	sub_wire1(82, 2)    <= sub_wire46(2);
	sub_wire1(82, 3)    <= sub_wire46(3);
	sub_wire1(82, 4)    <= sub_wire46(4);
	sub_wire1(82, 5)    <= sub_wire46(5);
	sub_wire1(82, 6)    <= sub_wire46(6);
	sub_wire1(82, 7)    <= sub_wire46(7);
	sub_wire1(82, 8)    <= sub_wire46(8);
	sub_wire1(82, 9)    <= sub_wire46(9);
	sub_wire1(82, 10)    <= sub_wire46(10);
	sub_wire1(82, 11)    <= sub_wire46(11);
	sub_wire1(82, 12)    <= sub_wire46(12);
	sub_wire1(82, 13)    <= sub_wire46(13);
	sub_wire1(82, 14)    <= sub_wire46(14);
	sub_wire1(82, 15)    <= sub_wire46(15);
	sub_wire1(82, 16)    <= sub_wire46(16);
	sub_wire1(82, 17)    <= sub_wire46(17);
	sub_wire1(82, 18)    <= sub_wire46(18);
	sub_wire1(82, 19)    <= sub_wire46(19);
	sub_wire1(82, 20)    <= sub_wire46(20);
	sub_wire1(82, 21)    <= sub_wire46(21);
	sub_wire1(82, 22)    <= sub_wire46(22);
	sub_wire1(82, 23)    <= sub_wire46(23);
	sub_wire1(82, 24)    <= sub_wire46(24);
	sub_wire1(82, 25)    <= sub_wire46(25);
	sub_wire1(82, 26)    <= sub_wire46(26);
	sub_wire1(82, 27)    <= sub_wire46(27);
	sub_wire1(82, 28)    <= sub_wire46(28);
	sub_wire1(82, 29)    <= sub_wire46(29);
	sub_wire1(82, 30)    <= sub_wire46(30);
	sub_wire1(82, 31)    <= sub_wire46(31);
	sub_wire1(81, 0)    <= sub_wire47(0);
	sub_wire1(81, 1)    <= sub_wire47(1);
	sub_wire1(81, 2)    <= sub_wire47(2);
	sub_wire1(81, 3)    <= sub_wire47(3);
	sub_wire1(81, 4)    <= sub_wire47(4);
	sub_wire1(81, 5)    <= sub_wire47(5);
	sub_wire1(81, 6)    <= sub_wire47(6);
	sub_wire1(81, 7)    <= sub_wire47(7);
	sub_wire1(81, 8)    <= sub_wire47(8);
	sub_wire1(81, 9)    <= sub_wire47(9);
	sub_wire1(81, 10)    <= sub_wire47(10);
	sub_wire1(81, 11)    <= sub_wire47(11);
	sub_wire1(81, 12)    <= sub_wire47(12);
	sub_wire1(81, 13)    <= sub_wire47(13);
	sub_wire1(81, 14)    <= sub_wire47(14);
	sub_wire1(81, 15)    <= sub_wire47(15);
	sub_wire1(81, 16)    <= sub_wire47(16);
	sub_wire1(81, 17)    <= sub_wire47(17);
	sub_wire1(81, 18)    <= sub_wire47(18);
	sub_wire1(81, 19)    <= sub_wire47(19);
	sub_wire1(81, 20)    <= sub_wire47(20);
	sub_wire1(81, 21)    <= sub_wire47(21);
	sub_wire1(81, 22)    <= sub_wire47(22);
	sub_wire1(81, 23)    <= sub_wire47(23);
	sub_wire1(81, 24)    <= sub_wire47(24);
	sub_wire1(81, 25)    <= sub_wire47(25);
	sub_wire1(81, 26)    <= sub_wire47(26);
	sub_wire1(81, 27)    <= sub_wire47(27);
	sub_wire1(81, 28)    <= sub_wire47(28);
	sub_wire1(81, 29)    <= sub_wire47(29);
	sub_wire1(81, 30)    <= sub_wire47(30);
	sub_wire1(81, 31)    <= sub_wire47(31);
	sub_wire1(80, 0)    <= sub_wire48(0);
	sub_wire1(80, 1)    <= sub_wire48(1);
	sub_wire1(80, 2)    <= sub_wire48(2);
	sub_wire1(80, 3)    <= sub_wire48(3);
	sub_wire1(80, 4)    <= sub_wire48(4);
	sub_wire1(80, 5)    <= sub_wire48(5);
	sub_wire1(80, 6)    <= sub_wire48(6);
	sub_wire1(80, 7)    <= sub_wire48(7);
	sub_wire1(80, 8)    <= sub_wire48(8);
	sub_wire1(80, 9)    <= sub_wire48(9);
	sub_wire1(80, 10)    <= sub_wire48(10);
	sub_wire1(80, 11)    <= sub_wire48(11);
	sub_wire1(80, 12)    <= sub_wire48(12);
	sub_wire1(80, 13)    <= sub_wire48(13);
	sub_wire1(80, 14)    <= sub_wire48(14);
	sub_wire1(80, 15)    <= sub_wire48(15);
	sub_wire1(80, 16)    <= sub_wire48(16);
	sub_wire1(80, 17)    <= sub_wire48(17);
	sub_wire1(80, 18)    <= sub_wire48(18);
	sub_wire1(80, 19)    <= sub_wire48(19);
	sub_wire1(80, 20)    <= sub_wire48(20);
	sub_wire1(80, 21)    <= sub_wire48(21);
	sub_wire1(80, 22)    <= sub_wire48(22);
	sub_wire1(80, 23)    <= sub_wire48(23);
	sub_wire1(80, 24)    <= sub_wire48(24);
	sub_wire1(80, 25)    <= sub_wire48(25);
	sub_wire1(80, 26)    <= sub_wire48(26);
	sub_wire1(80, 27)    <= sub_wire48(27);
	sub_wire1(80, 28)    <= sub_wire48(28);
	sub_wire1(80, 29)    <= sub_wire48(29);
	sub_wire1(80, 30)    <= sub_wire48(30);
	sub_wire1(80, 31)    <= sub_wire48(31);
	sub_wire1(79, 0)    <= sub_wire49(0);
	sub_wire1(79, 1)    <= sub_wire49(1);
	sub_wire1(79, 2)    <= sub_wire49(2);
	sub_wire1(79, 3)    <= sub_wire49(3);
	sub_wire1(79, 4)    <= sub_wire49(4);
	sub_wire1(79, 5)    <= sub_wire49(5);
	sub_wire1(79, 6)    <= sub_wire49(6);
	sub_wire1(79, 7)    <= sub_wire49(7);
	sub_wire1(79, 8)    <= sub_wire49(8);
	sub_wire1(79, 9)    <= sub_wire49(9);
	sub_wire1(79, 10)    <= sub_wire49(10);
	sub_wire1(79, 11)    <= sub_wire49(11);
	sub_wire1(79, 12)    <= sub_wire49(12);
	sub_wire1(79, 13)    <= sub_wire49(13);
	sub_wire1(79, 14)    <= sub_wire49(14);
	sub_wire1(79, 15)    <= sub_wire49(15);
	sub_wire1(79, 16)    <= sub_wire49(16);
	sub_wire1(79, 17)    <= sub_wire49(17);
	sub_wire1(79, 18)    <= sub_wire49(18);
	sub_wire1(79, 19)    <= sub_wire49(19);
	sub_wire1(79, 20)    <= sub_wire49(20);
	sub_wire1(79, 21)    <= sub_wire49(21);
	sub_wire1(79, 22)    <= sub_wire49(22);
	sub_wire1(79, 23)    <= sub_wire49(23);
	sub_wire1(79, 24)    <= sub_wire49(24);
	sub_wire1(79, 25)    <= sub_wire49(25);
	sub_wire1(79, 26)    <= sub_wire49(26);
	sub_wire1(79, 27)    <= sub_wire49(27);
	sub_wire1(79, 28)    <= sub_wire49(28);
	sub_wire1(79, 29)    <= sub_wire49(29);
	sub_wire1(79, 30)    <= sub_wire49(30);
	sub_wire1(79, 31)    <= sub_wire49(31);
	sub_wire1(78, 0)    <= sub_wire50(0);
	sub_wire1(78, 1)    <= sub_wire50(1);
	sub_wire1(78, 2)    <= sub_wire50(2);
	sub_wire1(78, 3)    <= sub_wire50(3);
	sub_wire1(78, 4)    <= sub_wire50(4);
	sub_wire1(78, 5)    <= sub_wire50(5);
	sub_wire1(78, 6)    <= sub_wire50(6);
	sub_wire1(78, 7)    <= sub_wire50(7);
	sub_wire1(78, 8)    <= sub_wire50(8);
	sub_wire1(78, 9)    <= sub_wire50(9);
	sub_wire1(78, 10)    <= sub_wire50(10);
	sub_wire1(78, 11)    <= sub_wire50(11);
	sub_wire1(78, 12)    <= sub_wire50(12);
	sub_wire1(78, 13)    <= sub_wire50(13);
	sub_wire1(78, 14)    <= sub_wire50(14);
	sub_wire1(78, 15)    <= sub_wire50(15);
	sub_wire1(78, 16)    <= sub_wire50(16);
	sub_wire1(78, 17)    <= sub_wire50(17);
	sub_wire1(78, 18)    <= sub_wire50(18);
	sub_wire1(78, 19)    <= sub_wire50(19);
	sub_wire1(78, 20)    <= sub_wire50(20);
	sub_wire1(78, 21)    <= sub_wire50(21);
	sub_wire1(78, 22)    <= sub_wire50(22);
	sub_wire1(78, 23)    <= sub_wire50(23);
	sub_wire1(78, 24)    <= sub_wire50(24);
	sub_wire1(78, 25)    <= sub_wire50(25);
	sub_wire1(78, 26)    <= sub_wire50(26);
	sub_wire1(78, 27)    <= sub_wire50(27);
	sub_wire1(78, 28)    <= sub_wire50(28);
	sub_wire1(78, 29)    <= sub_wire50(29);
	sub_wire1(78, 30)    <= sub_wire50(30);
	sub_wire1(78, 31)    <= sub_wire50(31);
	sub_wire1(77, 0)    <= sub_wire51(0);
	sub_wire1(77, 1)    <= sub_wire51(1);
	sub_wire1(77, 2)    <= sub_wire51(2);
	sub_wire1(77, 3)    <= sub_wire51(3);
	sub_wire1(77, 4)    <= sub_wire51(4);
	sub_wire1(77, 5)    <= sub_wire51(5);
	sub_wire1(77, 6)    <= sub_wire51(6);
	sub_wire1(77, 7)    <= sub_wire51(7);
	sub_wire1(77, 8)    <= sub_wire51(8);
	sub_wire1(77, 9)    <= sub_wire51(9);
	sub_wire1(77, 10)    <= sub_wire51(10);
	sub_wire1(77, 11)    <= sub_wire51(11);
	sub_wire1(77, 12)    <= sub_wire51(12);
	sub_wire1(77, 13)    <= sub_wire51(13);
	sub_wire1(77, 14)    <= sub_wire51(14);
	sub_wire1(77, 15)    <= sub_wire51(15);
	sub_wire1(77, 16)    <= sub_wire51(16);
	sub_wire1(77, 17)    <= sub_wire51(17);
	sub_wire1(77, 18)    <= sub_wire51(18);
	sub_wire1(77, 19)    <= sub_wire51(19);
	sub_wire1(77, 20)    <= sub_wire51(20);
	sub_wire1(77, 21)    <= sub_wire51(21);
	sub_wire1(77, 22)    <= sub_wire51(22);
	sub_wire1(77, 23)    <= sub_wire51(23);
	sub_wire1(77, 24)    <= sub_wire51(24);
	sub_wire1(77, 25)    <= sub_wire51(25);
	sub_wire1(77, 26)    <= sub_wire51(26);
	sub_wire1(77, 27)    <= sub_wire51(27);
	sub_wire1(77, 28)    <= sub_wire51(28);
	sub_wire1(77, 29)    <= sub_wire51(29);
	sub_wire1(77, 30)    <= sub_wire51(30);
	sub_wire1(77, 31)    <= sub_wire51(31);
	sub_wire1(76, 0)    <= sub_wire52(0);
	sub_wire1(76, 1)    <= sub_wire52(1);
	sub_wire1(76, 2)    <= sub_wire52(2);
	sub_wire1(76, 3)    <= sub_wire52(3);
	sub_wire1(76, 4)    <= sub_wire52(4);
	sub_wire1(76, 5)    <= sub_wire52(5);
	sub_wire1(76, 6)    <= sub_wire52(6);
	sub_wire1(76, 7)    <= sub_wire52(7);
	sub_wire1(76, 8)    <= sub_wire52(8);
	sub_wire1(76, 9)    <= sub_wire52(9);
	sub_wire1(76, 10)    <= sub_wire52(10);
	sub_wire1(76, 11)    <= sub_wire52(11);
	sub_wire1(76, 12)    <= sub_wire52(12);
	sub_wire1(76, 13)    <= sub_wire52(13);
	sub_wire1(76, 14)    <= sub_wire52(14);
	sub_wire1(76, 15)    <= sub_wire52(15);
	sub_wire1(76, 16)    <= sub_wire52(16);
	sub_wire1(76, 17)    <= sub_wire52(17);
	sub_wire1(76, 18)    <= sub_wire52(18);
	sub_wire1(76, 19)    <= sub_wire52(19);
	sub_wire1(76, 20)    <= sub_wire52(20);
	sub_wire1(76, 21)    <= sub_wire52(21);
	sub_wire1(76, 22)    <= sub_wire52(22);
	sub_wire1(76, 23)    <= sub_wire52(23);
	sub_wire1(76, 24)    <= sub_wire52(24);
	sub_wire1(76, 25)    <= sub_wire52(25);
	sub_wire1(76, 26)    <= sub_wire52(26);
	sub_wire1(76, 27)    <= sub_wire52(27);
	sub_wire1(76, 28)    <= sub_wire52(28);
	sub_wire1(76, 29)    <= sub_wire52(29);
	sub_wire1(76, 30)    <= sub_wire52(30);
	sub_wire1(76, 31)    <= sub_wire52(31);
	sub_wire1(75, 0)    <= sub_wire53(0);
	sub_wire1(75, 1)    <= sub_wire53(1);
	sub_wire1(75, 2)    <= sub_wire53(2);
	sub_wire1(75, 3)    <= sub_wire53(3);
	sub_wire1(75, 4)    <= sub_wire53(4);
	sub_wire1(75, 5)    <= sub_wire53(5);
	sub_wire1(75, 6)    <= sub_wire53(6);
	sub_wire1(75, 7)    <= sub_wire53(7);
	sub_wire1(75, 8)    <= sub_wire53(8);
	sub_wire1(75, 9)    <= sub_wire53(9);
	sub_wire1(75, 10)    <= sub_wire53(10);
	sub_wire1(75, 11)    <= sub_wire53(11);
	sub_wire1(75, 12)    <= sub_wire53(12);
	sub_wire1(75, 13)    <= sub_wire53(13);
	sub_wire1(75, 14)    <= sub_wire53(14);
	sub_wire1(75, 15)    <= sub_wire53(15);
	sub_wire1(75, 16)    <= sub_wire53(16);
	sub_wire1(75, 17)    <= sub_wire53(17);
	sub_wire1(75, 18)    <= sub_wire53(18);
	sub_wire1(75, 19)    <= sub_wire53(19);
	sub_wire1(75, 20)    <= sub_wire53(20);
	sub_wire1(75, 21)    <= sub_wire53(21);
	sub_wire1(75, 22)    <= sub_wire53(22);
	sub_wire1(75, 23)    <= sub_wire53(23);
	sub_wire1(75, 24)    <= sub_wire53(24);
	sub_wire1(75, 25)    <= sub_wire53(25);
	sub_wire1(75, 26)    <= sub_wire53(26);
	sub_wire1(75, 27)    <= sub_wire53(27);
	sub_wire1(75, 28)    <= sub_wire53(28);
	sub_wire1(75, 29)    <= sub_wire53(29);
	sub_wire1(75, 30)    <= sub_wire53(30);
	sub_wire1(75, 31)    <= sub_wire53(31);
	sub_wire1(74, 0)    <= sub_wire54(0);
	sub_wire1(74, 1)    <= sub_wire54(1);
	sub_wire1(74, 2)    <= sub_wire54(2);
	sub_wire1(74, 3)    <= sub_wire54(3);
	sub_wire1(74, 4)    <= sub_wire54(4);
	sub_wire1(74, 5)    <= sub_wire54(5);
	sub_wire1(74, 6)    <= sub_wire54(6);
	sub_wire1(74, 7)    <= sub_wire54(7);
	sub_wire1(74, 8)    <= sub_wire54(8);
	sub_wire1(74, 9)    <= sub_wire54(9);
	sub_wire1(74, 10)    <= sub_wire54(10);
	sub_wire1(74, 11)    <= sub_wire54(11);
	sub_wire1(74, 12)    <= sub_wire54(12);
	sub_wire1(74, 13)    <= sub_wire54(13);
	sub_wire1(74, 14)    <= sub_wire54(14);
	sub_wire1(74, 15)    <= sub_wire54(15);
	sub_wire1(74, 16)    <= sub_wire54(16);
	sub_wire1(74, 17)    <= sub_wire54(17);
	sub_wire1(74, 18)    <= sub_wire54(18);
	sub_wire1(74, 19)    <= sub_wire54(19);
	sub_wire1(74, 20)    <= sub_wire54(20);
	sub_wire1(74, 21)    <= sub_wire54(21);
	sub_wire1(74, 22)    <= sub_wire54(22);
	sub_wire1(74, 23)    <= sub_wire54(23);
	sub_wire1(74, 24)    <= sub_wire54(24);
	sub_wire1(74, 25)    <= sub_wire54(25);
	sub_wire1(74, 26)    <= sub_wire54(26);
	sub_wire1(74, 27)    <= sub_wire54(27);
	sub_wire1(74, 28)    <= sub_wire54(28);
	sub_wire1(74, 29)    <= sub_wire54(29);
	sub_wire1(74, 30)    <= sub_wire54(30);
	sub_wire1(74, 31)    <= sub_wire54(31);
	sub_wire1(73, 0)    <= sub_wire55(0);
	sub_wire1(73, 1)    <= sub_wire55(1);
	sub_wire1(73, 2)    <= sub_wire55(2);
	sub_wire1(73, 3)    <= sub_wire55(3);
	sub_wire1(73, 4)    <= sub_wire55(4);
	sub_wire1(73, 5)    <= sub_wire55(5);
	sub_wire1(73, 6)    <= sub_wire55(6);
	sub_wire1(73, 7)    <= sub_wire55(7);
	sub_wire1(73, 8)    <= sub_wire55(8);
	sub_wire1(73, 9)    <= sub_wire55(9);
	sub_wire1(73, 10)    <= sub_wire55(10);
	sub_wire1(73, 11)    <= sub_wire55(11);
	sub_wire1(73, 12)    <= sub_wire55(12);
	sub_wire1(73, 13)    <= sub_wire55(13);
	sub_wire1(73, 14)    <= sub_wire55(14);
	sub_wire1(73, 15)    <= sub_wire55(15);
	sub_wire1(73, 16)    <= sub_wire55(16);
	sub_wire1(73, 17)    <= sub_wire55(17);
	sub_wire1(73, 18)    <= sub_wire55(18);
	sub_wire1(73, 19)    <= sub_wire55(19);
	sub_wire1(73, 20)    <= sub_wire55(20);
	sub_wire1(73, 21)    <= sub_wire55(21);
	sub_wire1(73, 22)    <= sub_wire55(22);
	sub_wire1(73, 23)    <= sub_wire55(23);
	sub_wire1(73, 24)    <= sub_wire55(24);
	sub_wire1(73, 25)    <= sub_wire55(25);
	sub_wire1(73, 26)    <= sub_wire55(26);
	sub_wire1(73, 27)    <= sub_wire55(27);
	sub_wire1(73, 28)    <= sub_wire55(28);
	sub_wire1(73, 29)    <= sub_wire55(29);
	sub_wire1(73, 30)    <= sub_wire55(30);
	sub_wire1(73, 31)    <= sub_wire55(31);
	sub_wire1(72, 0)    <= sub_wire56(0);
	sub_wire1(72, 1)    <= sub_wire56(1);
	sub_wire1(72, 2)    <= sub_wire56(2);
	sub_wire1(72, 3)    <= sub_wire56(3);
	sub_wire1(72, 4)    <= sub_wire56(4);
	sub_wire1(72, 5)    <= sub_wire56(5);
	sub_wire1(72, 6)    <= sub_wire56(6);
	sub_wire1(72, 7)    <= sub_wire56(7);
	sub_wire1(72, 8)    <= sub_wire56(8);
	sub_wire1(72, 9)    <= sub_wire56(9);
	sub_wire1(72, 10)    <= sub_wire56(10);
	sub_wire1(72, 11)    <= sub_wire56(11);
	sub_wire1(72, 12)    <= sub_wire56(12);
	sub_wire1(72, 13)    <= sub_wire56(13);
	sub_wire1(72, 14)    <= sub_wire56(14);
	sub_wire1(72, 15)    <= sub_wire56(15);
	sub_wire1(72, 16)    <= sub_wire56(16);
	sub_wire1(72, 17)    <= sub_wire56(17);
	sub_wire1(72, 18)    <= sub_wire56(18);
	sub_wire1(72, 19)    <= sub_wire56(19);
	sub_wire1(72, 20)    <= sub_wire56(20);
	sub_wire1(72, 21)    <= sub_wire56(21);
	sub_wire1(72, 22)    <= sub_wire56(22);
	sub_wire1(72, 23)    <= sub_wire56(23);
	sub_wire1(72, 24)    <= sub_wire56(24);
	sub_wire1(72, 25)    <= sub_wire56(25);
	sub_wire1(72, 26)    <= sub_wire56(26);
	sub_wire1(72, 27)    <= sub_wire56(27);
	sub_wire1(72, 28)    <= sub_wire56(28);
	sub_wire1(72, 29)    <= sub_wire56(29);
	sub_wire1(72, 30)    <= sub_wire56(30);
	sub_wire1(72, 31)    <= sub_wire56(31);
	sub_wire1(71, 0)    <= sub_wire57(0);
	sub_wire1(71, 1)    <= sub_wire57(1);
	sub_wire1(71, 2)    <= sub_wire57(2);
	sub_wire1(71, 3)    <= sub_wire57(3);
	sub_wire1(71, 4)    <= sub_wire57(4);
	sub_wire1(71, 5)    <= sub_wire57(5);
	sub_wire1(71, 6)    <= sub_wire57(6);
	sub_wire1(71, 7)    <= sub_wire57(7);
	sub_wire1(71, 8)    <= sub_wire57(8);
	sub_wire1(71, 9)    <= sub_wire57(9);
	sub_wire1(71, 10)    <= sub_wire57(10);
	sub_wire1(71, 11)    <= sub_wire57(11);
	sub_wire1(71, 12)    <= sub_wire57(12);
	sub_wire1(71, 13)    <= sub_wire57(13);
	sub_wire1(71, 14)    <= sub_wire57(14);
	sub_wire1(71, 15)    <= sub_wire57(15);
	sub_wire1(71, 16)    <= sub_wire57(16);
	sub_wire1(71, 17)    <= sub_wire57(17);
	sub_wire1(71, 18)    <= sub_wire57(18);
	sub_wire1(71, 19)    <= sub_wire57(19);
	sub_wire1(71, 20)    <= sub_wire57(20);
	sub_wire1(71, 21)    <= sub_wire57(21);
	sub_wire1(71, 22)    <= sub_wire57(22);
	sub_wire1(71, 23)    <= sub_wire57(23);
	sub_wire1(71, 24)    <= sub_wire57(24);
	sub_wire1(71, 25)    <= sub_wire57(25);
	sub_wire1(71, 26)    <= sub_wire57(26);
	sub_wire1(71, 27)    <= sub_wire57(27);
	sub_wire1(71, 28)    <= sub_wire57(28);
	sub_wire1(71, 29)    <= sub_wire57(29);
	sub_wire1(71, 30)    <= sub_wire57(30);
	sub_wire1(71, 31)    <= sub_wire57(31);
	sub_wire1(70, 0)    <= sub_wire58(0);
	sub_wire1(70, 1)    <= sub_wire58(1);
	sub_wire1(70, 2)    <= sub_wire58(2);
	sub_wire1(70, 3)    <= sub_wire58(3);
	sub_wire1(70, 4)    <= sub_wire58(4);
	sub_wire1(70, 5)    <= sub_wire58(5);
	sub_wire1(70, 6)    <= sub_wire58(6);
	sub_wire1(70, 7)    <= sub_wire58(7);
	sub_wire1(70, 8)    <= sub_wire58(8);
	sub_wire1(70, 9)    <= sub_wire58(9);
	sub_wire1(70, 10)    <= sub_wire58(10);
	sub_wire1(70, 11)    <= sub_wire58(11);
	sub_wire1(70, 12)    <= sub_wire58(12);
	sub_wire1(70, 13)    <= sub_wire58(13);
	sub_wire1(70, 14)    <= sub_wire58(14);
	sub_wire1(70, 15)    <= sub_wire58(15);
	sub_wire1(70, 16)    <= sub_wire58(16);
	sub_wire1(70, 17)    <= sub_wire58(17);
	sub_wire1(70, 18)    <= sub_wire58(18);
	sub_wire1(70, 19)    <= sub_wire58(19);
	sub_wire1(70, 20)    <= sub_wire58(20);
	sub_wire1(70, 21)    <= sub_wire58(21);
	sub_wire1(70, 22)    <= sub_wire58(22);
	sub_wire1(70, 23)    <= sub_wire58(23);
	sub_wire1(70, 24)    <= sub_wire58(24);
	sub_wire1(70, 25)    <= sub_wire58(25);
	sub_wire1(70, 26)    <= sub_wire58(26);
	sub_wire1(70, 27)    <= sub_wire58(27);
	sub_wire1(70, 28)    <= sub_wire58(28);
	sub_wire1(70, 29)    <= sub_wire58(29);
	sub_wire1(70, 30)    <= sub_wire58(30);
	sub_wire1(70, 31)    <= sub_wire58(31);
	sub_wire1(69, 0)    <= sub_wire59(0);
	sub_wire1(69, 1)    <= sub_wire59(1);
	sub_wire1(69, 2)    <= sub_wire59(2);
	sub_wire1(69, 3)    <= sub_wire59(3);
	sub_wire1(69, 4)    <= sub_wire59(4);
	sub_wire1(69, 5)    <= sub_wire59(5);
	sub_wire1(69, 6)    <= sub_wire59(6);
	sub_wire1(69, 7)    <= sub_wire59(7);
	sub_wire1(69, 8)    <= sub_wire59(8);
	sub_wire1(69, 9)    <= sub_wire59(9);
	sub_wire1(69, 10)    <= sub_wire59(10);
	sub_wire1(69, 11)    <= sub_wire59(11);
	sub_wire1(69, 12)    <= sub_wire59(12);
	sub_wire1(69, 13)    <= sub_wire59(13);
	sub_wire1(69, 14)    <= sub_wire59(14);
	sub_wire1(69, 15)    <= sub_wire59(15);
	sub_wire1(69, 16)    <= sub_wire59(16);
	sub_wire1(69, 17)    <= sub_wire59(17);
	sub_wire1(69, 18)    <= sub_wire59(18);
	sub_wire1(69, 19)    <= sub_wire59(19);
	sub_wire1(69, 20)    <= sub_wire59(20);
	sub_wire1(69, 21)    <= sub_wire59(21);
	sub_wire1(69, 22)    <= sub_wire59(22);
	sub_wire1(69, 23)    <= sub_wire59(23);
	sub_wire1(69, 24)    <= sub_wire59(24);
	sub_wire1(69, 25)    <= sub_wire59(25);
	sub_wire1(69, 26)    <= sub_wire59(26);
	sub_wire1(69, 27)    <= sub_wire59(27);
	sub_wire1(69, 28)    <= sub_wire59(28);
	sub_wire1(69, 29)    <= sub_wire59(29);
	sub_wire1(69, 30)    <= sub_wire59(30);
	sub_wire1(69, 31)    <= sub_wire59(31);
	sub_wire1(68, 0)    <= sub_wire60(0);
	sub_wire1(68, 1)    <= sub_wire60(1);
	sub_wire1(68, 2)    <= sub_wire60(2);
	sub_wire1(68, 3)    <= sub_wire60(3);
	sub_wire1(68, 4)    <= sub_wire60(4);
	sub_wire1(68, 5)    <= sub_wire60(5);
	sub_wire1(68, 6)    <= sub_wire60(6);
	sub_wire1(68, 7)    <= sub_wire60(7);
	sub_wire1(68, 8)    <= sub_wire60(8);
	sub_wire1(68, 9)    <= sub_wire60(9);
	sub_wire1(68, 10)    <= sub_wire60(10);
	sub_wire1(68, 11)    <= sub_wire60(11);
	sub_wire1(68, 12)    <= sub_wire60(12);
	sub_wire1(68, 13)    <= sub_wire60(13);
	sub_wire1(68, 14)    <= sub_wire60(14);
	sub_wire1(68, 15)    <= sub_wire60(15);
	sub_wire1(68, 16)    <= sub_wire60(16);
	sub_wire1(68, 17)    <= sub_wire60(17);
	sub_wire1(68, 18)    <= sub_wire60(18);
	sub_wire1(68, 19)    <= sub_wire60(19);
	sub_wire1(68, 20)    <= sub_wire60(20);
	sub_wire1(68, 21)    <= sub_wire60(21);
	sub_wire1(68, 22)    <= sub_wire60(22);
	sub_wire1(68, 23)    <= sub_wire60(23);
	sub_wire1(68, 24)    <= sub_wire60(24);
	sub_wire1(68, 25)    <= sub_wire60(25);
	sub_wire1(68, 26)    <= sub_wire60(26);
	sub_wire1(68, 27)    <= sub_wire60(27);
	sub_wire1(68, 28)    <= sub_wire60(28);
	sub_wire1(68, 29)    <= sub_wire60(29);
	sub_wire1(68, 30)    <= sub_wire60(30);
	sub_wire1(68, 31)    <= sub_wire60(31);
	sub_wire1(67, 0)    <= sub_wire61(0);
	sub_wire1(67, 1)    <= sub_wire61(1);
	sub_wire1(67, 2)    <= sub_wire61(2);
	sub_wire1(67, 3)    <= sub_wire61(3);
	sub_wire1(67, 4)    <= sub_wire61(4);
	sub_wire1(67, 5)    <= sub_wire61(5);
	sub_wire1(67, 6)    <= sub_wire61(6);
	sub_wire1(67, 7)    <= sub_wire61(7);
	sub_wire1(67, 8)    <= sub_wire61(8);
	sub_wire1(67, 9)    <= sub_wire61(9);
	sub_wire1(67, 10)    <= sub_wire61(10);
	sub_wire1(67, 11)    <= sub_wire61(11);
	sub_wire1(67, 12)    <= sub_wire61(12);
	sub_wire1(67, 13)    <= sub_wire61(13);
	sub_wire1(67, 14)    <= sub_wire61(14);
	sub_wire1(67, 15)    <= sub_wire61(15);
	sub_wire1(67, 16)    <= sub_wire61(16);
	sub_wire1(67, 17)    <= sub_wire61(17);
	sub_wire1(67, 18)    <= sub_wire61(18);
	sub_wire1(67, 19)    <= sub_wire61(19);
	sub_wire1(67, 20)    <= sub_wire61(20);
	sub_wire1(67, 21)    <= sub_wire61(21);
	sub_wire1(67, 22)    <= sub_wire61(22);
	sub_wire1(67, 23)    <= sub_wire61(23);
	sub_wire1(67, 24)    <= sub_wire61(24);
	sub_wire1(67, 25)    <= sub_wire61(25);
	sub_wire1(67, 26)    <= sub_wire61(26);
	sub_wire1(67, 27)    <= sub_wire61(27);
	sub_wire1(67, 28)    <= sub_wire61(28);
	sub_wire1(67, 29)    <= sub_wire61(29);
	sub_wire1(67, 30)    <= sub_wire61(30);
	sub_wire1(67, 31)    <= sub_wire61(31);
	sub_wire1(66, 0)    <= sub_wire62(0);
	sub_wire1(66, 1)    <= sub_wire62(1);
	sub_wire1(66, 2)    <= sub_wire62(2);
	sub_wire1(66, 3)    <= sub_wire62(3);
	sub_wire1(66, 4)    <= sub_wire62(4);
	sub_wire1(66, 5)    <= sub_wire62(5);
	sub_wire1(66, 6)    <= sub_wire62(6);
	sub_wire1(66, 7)    <= sub_wire62(7);
	sub_wire1(66, 8)    <= sub_wire62(8);
	sub_wire1(66, 9)    <= sub_wire62(9);
	sub_wire1(66, 10)    <= sub_wire62(10);
	sub_wire1(66, 11)    <= sub_wire62(11);
	sub_wire1(66, 12)    <= sub_wire62(12);
	sub_wire1(66, 13)    <= sub_wire62(13);
	sub_wire1(66, 14)    <= sub_wire62(14);
	sub_wire1(66, 15)    <= sub_wire62(15);
	sub_wire1(66, 16)    <= sub_wire62(16);
	sub_wire1(66, 17)    <= sub_wire62(17);
	sub_wire1(66, 18)    <= sub_wire62(18);
	sub_wire1(66, 19)    <= sub_wire62(19);
	sub_wire1(66, 20)    <= sub_wire62(20);
	sub_wire1(66, 21)    <= sub_wire62(21);
	sub_wire1(66, 22)    <= sub_wire62(22);
	sub_wire1(66, 23)    <= sub_wire62(23);
	sub_wire1(66, 24)    <= sub_wire62(24);
	sub_wire1(66, 25)    <= sub_wire62(25);
	sub_wire1(66, 26)    <= sub_wire62(26);
	sub_wire1(66, 27)    <= sub_wire62(27);
	sub_wire1(66, 28)    <= sub_wire62(28);
	sub_wire1(66, 29)    <= sub_wire62(29);
	sub_wire1(66, 30)    <= sub_wire62(30);
	sub_wire1(66, 31)    <= sub_wire62(31);
	sub_wire1(65, 0)    <= sub_wire63(0);
	sub_wire1(65, 1)    <= sub_wire63(1);
	sub_wire1(65, 2)    <= sub_wire63(2);
	sub_wire1(65, 3)    <= sub_wire63(3);
	sub_wire1(65, 4)    <= sub_wire63(4);
	sub_wire1(65, 5)    <= sub_wire63(5);
	sub_wire1(65, 6)    <= sub_wire63(6);
	sub_wire1(65, 7)    <= sub_wire63(7);
	sub_wire1(65, 8)    <= sub_wire63(8);
	sub_wire1(65, 9)    <= sub_wire63(9);
	sub_wire1(65, 10)    <= sub_wire63(10);
	sub_wire1(65, 11)    <= sub_wire63(11);
	sub_wire1(65, 12)    <= sub_wire63(12);
	sub_wire1(65, 13)    <= sub_wire63(13);
	sub_wire1(65, 14)    <= sub_wire63(14);
	sub_wire1(65, 15)    <= sub_wire63(15);
	sub_wire1(65, 16)    <= sub_wire63(16);
	sub_wire1(65, 17)    <= sub_wire63(17);
	sub_wire1(65, 18)    <= sub_wire63(18);
	sub_wire1(65, 19)    <= sub_wire63(19);
	sub_wire1(65, 20)    <= sub_wire63(20);
	sub_wire1(65, 21)    <= sub_wire63(21);
	sub_wire1(65, 22)    <= sub_wire63(22);
	sub_wire1(65, 23)    <= sub_wire63(23);
	sub_wire1(65, 24)    <= sub_wire63(24);
	sub_wire1(65, 25)    <= sub_wire63(25);
	sub_wire1(65, 26)    <= sub_wire63(26);
	sub_wire1(65, 27)    <= sub_wire63(27);
	sub_wire1(65, 28)    <= sub_wire63(28);
	sub_wire1(65, 29)    <= sub_wire63(29);
	sub_wire1(65, 30)    <= sub_wire63(30);
	sub_wire1(65, 31)    <= sub_wire63(31);
	sub_wire1(64, 0)    <= sub_wire64(0);
	sub_wire1(64, 1)    <= sub_wire64(1);
	sub_wire1(64, 2)    <= sub_wire64(2);
	sub_wire1(64, 3)    <= sub_wire64(3);
	sub_wire1(64, 4)    <= sub_wire64(4);
	sub_wire1(64, 5)    <= sub_wire64(5);
	sub_wire1(64, 6)    <= sub_wire64(6);
	sub_wire1(64, 7)    <= sub_wire64(7);
	sub_wire1(64, 8)    <= sub_wire64(8);
	sub_wire1(64, 9)    <= sub_wire64(9);
	sub_wire1(64, 10)    <= sub_wire64(10);
	sub_wire1(64, 11)    <= sub_wire64(11);
	sub_wire1(64, 12)    <= sub_wire64(12);
	sub_wire1(64, 13)    <= sub_wire64(13);
	sub_wire1(64, 14)    <= sub_wire64(14);
	sub_wire1(64, 15)    <= sub_wire64(15);
	sub_wire1(64, 16)    <= sub_wire64(16);
	sub_wire1(64, 17)    <= sub_wire64(17);
	sub_wire1(64, 18)    <= sub_wire64(18);
	sub_wire1(64, 19)    <= sub_wire64(19);
	sub_wire1(64, 20)    <= sub_wire64(20);
	sub_wire1(64, 21)    <= sub_wire64(21);
	sub_wire1(64, 22)    <= sub_wire64(22);
	sub_wire1(64, 23)    <= sub_wire64(23);
	sub_wire1(64, 24)    <= sub_wire64(24);
	sub_wire1(64, 25)    <= sub_wire64(25);
	sub_wire1(64, 26)    <= sub_wire64(26);
	sub_wire1(64, 27)    <= sub_wire64(27);
	sub_wire1(64, 28)    <= sub_wire64(28);
	sub_wire1(64, 29)    <= sub_wire64(29);
	sub_wire1(64, 30)    <= sub_wire64(30);
	sub_wire1(64, 31)    <= sub_wire64(31);
	sub_wire1(63, 0)    <= sub_wire65(0);
	sub_wire1(63, 1)    <= sub_wire65(1);
	sub_wire1(63, 2)    <= sub_wire65(2);
	sub_wire1(63, 3)    <= sub_wire65(3);
	sub_wire1(63, 4)    <= sub_wire65(4);
	sub_wire1(63, 5)    <= sub_wire65(5);
	sub_wire1(63, 6)    <= sub_wire65(6);
	sub_wire1(63, 7)    <= sub_wire65(7);
	sub_wire1(63, 8)    <= sub_wire65(8);
	sub_wire1(63, 9)    <= sub_wire65(9);
	sub_wire1(63, 10)    <= sub_wire65(10);
	sub_wire1(63, 11)    <= sub_wire65(11);
	sub_wire1(63, 12)    <= sub_wire65(12);
	sub_wire1(63, 13)    <= sub_wire65(13);
	sub_wire1(63, 14)    <= sub_wire65(14);
	sub_wire1(63, 15)    <= sub_wire65(15);
	sub_wire1(63, 16)    <= sub_wire65(16);
	sub_wire1(63, 17)    <= sub_wire65(17);
	sub_wire1(63, 18)    <= sub_wire65(18);
	sub_wire1(63, 19)    <= sub_wire65(19);
	sub_wire1(63, 20)    <= sub_wire65(20);
	sub_wire1(63, 21)    <= sub_wire65(21);
	sub_wire1(63, 22)    <= sub_wire65(22);
	sub_wire1(63, 23)    <= sub_wire65(23);
	sub_wire1(63, 24)    <= sub_wire65(24);
	sub_wire1(63, 25)    <= sub_wire65(25);
	sub_wire1(63, 26)    <= sub_wire65(26);
	sub_wire1(63, 27)    <= sub_wire65(27);
	sub_wire1(63, 28)    <= sub_wire65(28);
	sub_wire1(63, 29)    <= sub_wire65(29);
	sub_wire1(63, 30)    <= sub_wire65(30);
	sub_wire1(63, 31)    <= sub_wire65(31);
	sub_wire1(62, 0)    <= sub_wire66(0);
	sub_wire1(62, 1)    <= sub_wire66(1);
	sub_wire1(62, 2)    <= sub_wire66(2);
	sub_wire1(62, 3)    <= sub_wire66(3);
	sub_wire1(62, 4)    <= sub_wire66(4);
	sub_wire1(62, 5)    <= sub_wire66(5);
	sub_wire1(62, 6)    <= sub_wire66(6);
	sub_wire1(62, 7)    <= sub_wire66(7);
	sub_wire1(62, 8)    <= sub_wire66(8);
	sub_wire1(62, 9)    <= sub_wire66(9);
	sub_wire1(62, 10)    <= sub_wire66(10);
	sub_wire1(62, 11)    <= sub_wire66(11);
	sub_wire1(62, 12)    <= sub_wire66(12);
	sub_wire1(62, 13)    <= sub_wire66(13);
	sub_wire1(62, 14)    <= sub_wire66(14);
	sub_wire1(62, 15)    <= sub_wire66(15);
	sub_wire1(62, 16)    <= sub_wire66(16);
	sub_wire1(62, 17)    <= sub_wire66(17);
	sub_wire1(62, 18)    <= sub_wire66(18);
	sub_wire1(62, 19)    <= sub_wire66(19);
	sub_wire1(62, 20)    <= sub_wire66(20);
	sub_wire1(62, 21)    <= sub_wire66(21);
	sub_wire1(62, 22)    <= sub_wire66(22);
	sub_wire1(62, 23)    <= sub_wire66(23);
	sub_wire1(62, 24)    <= sub_wire66(24);
	sub_wire1(62, 25)    <= sub_wire66(25);
	sub_wire1(62, 26)    <= sub_wire66(26);
	sub_wire1(62, 27)    <= sub_wire66(27);
	sub_wire1(62, 28)    <= sub_wire66(28);
	sub_wire1(62, 29)    <= sub_wire66(29);
	sub_wire1(62, 30)    <= sub_wire66(30);
	sub_wire1(62, 31)    <= sub_wire66(31);
	sub_wire1(61, 0)    <= sub_wire67(0);
	sub_wire1(61, 1)    <= sub_wire67(1);
	sub_wire1(61, 2)    <= sub_wire67(2);
	sub_wire1(61, 3)    <= sub_wire67(3);
	sub_wire1(61, 4)    <= sub_wire67(4);
	sub_wire1(61, 5)    <= sub_wire67(5);
	sub_wire1(61, 6)    <= sub_wire67(6);
	sub_wire1(61, 7)    <= sub_wire67(7);
	sub_wire1(61, 8)    <= sub_wire67(8);
	sub_wire1(61, 9)    <= sub_wire67(9);
	sub_wire1(61, 10)    <= sub_wire67(10);
	sub_wire1(61, 11)    <= sub_wire67(11);
	sub_wire1(61, 12)    <= sub_wire67(12);
	sub_wire1(61, 13)    <= sub_wire67(13);
	sub_wire1(61, 14)    <= sub_wire67(14);
	sub_wire1(61, 15)    <= sub_wire67(15);
	sub_wire1(61, 16)    <= sub_wire67(16);
	sub_wire1(61, 17)    <= sub_wire67(17);
	sub_wire1(61, 18)    <= sub_wire67(18);
	sub_wire1(61, 19)    <= sub_wire67(19);
	sub_wire1(61, 20)    <= sub_wire67(20);
	sub_wire1(61, 21)    <= sub_wire67(21);
	sub_wire1(61, 22)    <= sub_wire67(22);
	sub_wire1(61, 23)    <= sub_wire67(23);
	sub_wire1(61, 24)    <= sub_wire67(24);
	sub_wire1(61, 25)    <= sub_wire67(25);
	sub_wire1(61, 26)    <= sub_wire67(26);
	sub_wire1(61, 27)    <= sub_wire67(27);
	sub_wire1(61, 28)    <= sub_wire67(28);
	sub_wire1(61, 29)    <= sub_wire67(29);
	sub_wire1(61, 30)    <= sub_wire67(30);
	sub_wire1(61, 31)    <= sub_wire67(31);
	sub_wire1(60, 0)    <= sub_wire68(0);
	sub_wire1(60, 1)    <= sub_wire68(1);
	sub_wire1(60, 2)    <= sub_wire68(2);
	sub_wire1(60, 3)    <= sub_wire68(3);
	sub_wire1(60, 4)    <= sub_wire68(4);
	sub_wire1(60, 5)    <= sub_wire68(5);
	sub_wire1(60, 6)    <= sub_wire68(6);
	sub_wire1(60, 7)    <= sub_wire68(7);
	sub_wire1(60, 8)    <= sub_wire68(8);
	sub_wire1(60, 9)    <= sub_wire68(9);
	sub_wire1(60, 10)    <= sub_wire68(10);
	sub_wire1(60, 11)    <= sub_wire68(11);
	sub_wire1(60, 12)    <= sub_wire68(12);
	sub_wire1(60, 13)    <= sub_wire68(13);
	sub_wire1(60, 14)    <= sub_wire68(14);
	sub_wire1(60, 15)    <= sub_wire68(15);
	sub_wire1(60, 16)    <= sub_wire68(16);
	sub_wire1(60, 17)    <= sub_wire68(17);
	sub_wire1(60, 18)    <= sub_wire68(18);
	sub_wire1(60, 19)    <= sub_wire68(19);
	sub_wire1(60, 20)    <= sub_wire68(20);
	sub_wire1(60, 21)    <= sub_wire68(21);
	sub_wire1(60, 22)    <= sub_wire68(22);
	sub_wire1(60, 23)    <= sub_wire68(23);
	sub_wire1(60, 24)    <= sub_wire68(24);
	sub_wire1(60, 25)    <= sub_wire68(25);
	sub_wire1(60, 26)    <= sub_wire68(26);
	sub_wire1(60, 27)    <= sub_wire68(27);
	sub_wire1(60, 28)    <= sub_wire68(28);
	sub_wire1(60, 29)    <= sub_wire68(29);
	sub_wire1(60, 30)    <= sub_wire68(30);
	sub_wire1(60, 31)    <= sub_wire68(31);
	sub_wire1(59, 0)    <= sub_wire69(0);
	sub_wire1(59, 1)    <= sub_wire69(1);
	sub_wire1(59, 2)    <= sub_wire69(2);
	sub_wire1(59, 3)    <= sub_wire69(3);
	sub_wire1(59, 4)    <= sub_wire69(4);
	sub_wire1(59, 5)    <= sub_wire69(5);
	sub_wire1(59, 6)    <= sub_wire69(6);
	sub_wire1(59, 7)    <= sub_wire69(7);
	sub_wire1(59, 8)    <= sub_wire69(8);
	sub_wire1(59, 9)    <= sub_wire69(9);
	sub_wire1(59, 10)    <= sub_wire69(10);
	sub_wire1(59, 11)    <= sub_wire69(11);
	sub_wire1(59, 12)    <= sub_wire69(12);
	sub_wire1(59, 13)    <= sub_wire69(13);
	sub_wire1(59, 14)    <= sub_wire69(14);
	sub_wire1(59, 15)    <= sub_wire69(15);
	sub_wire1(59, 16)    <= sub_wire69(16);
	sub_wire1(59, 17)    <= sub_wire69(17);
	sub_wire1(59, 18)    <= sub_wire69(18);
	sub_wire1(59, 19)    <= sub_wire69(19);
	sub_wire1(59, 20)    <= sub_wire69(20);
	sub_wire1(59, 21)    <= sub_wire69(21);
	sub_wire1(59, 22)    <= sub_wire69(22);
	sub_wire1(59, 23)    <= sub_wire69(23);
	sub_wire1(59, 24)    <= sub_wire69(24);
	sub_wire1(59, 25)    <= sub_wire69(25);
	sub_wire1(59, 26)    <= sub_wire69(26);
	sub_wire1(59, 27)    <= sub_wire69(27);
	sub_wire1(59, 28)    <= sub_wire69(28);
	sub_wire1(59, 29)    <= sub_wire69(29);
	sub_wire1(59, 30)    <= sub_wire69(30);
	sub_wire1(59, 31)    <= sub_wire69(31);
	sub_wire1(58, 0)    <= sub_wire70(0);
	sub_wire1(58, 1)    <= sub_wire70(1);
	sub_wire1(58, 2)    <= sub_wire70(2);
	sub_wire1(58, 3)    <= sub_wire70(3);
	sub_wire1(58, 4)    <= sub_wire70(4);
	sub_wire1(58, 5)    <= sub_wire70(5);
	sub_wire1(58, 6)    <= sub_wire70(6);
	sub_wire1(58, 7)    <= sub_wire70(7);
	sub_wire1(58, 8)    <= sub_wire70(8);
	sub_wire1(58, 9)    <= sub_wire70(9);
	sub_wire1(58, 10)    <= sub_wire70(10);
	sub_wire1(58, 11)    <= sub_wire70(11);
	sub_wire1(58, 12)    <= sub_wire70(12);
	sub_wire1(58, 13)    <= sub_wire70(13);
	sub_wire1(58, 14)    <= sub_wire70(14);
	sub_wire1(58, 15)    <= sub_wire70(15);
	sub_wire1(58, 16)    <= sub_wire70(16);
	sub_wire1(58, 17)    <= sub_wire70(17);
	sub_wire1(58, 18)    <= sub_wire70(18);
	sub_wire1(58, 19)    <= sub_wire70(19);
	sub_wire1(58, 20)    <= sub_wire70(20);
	sub_wire1(58, 21)    <= sub_wire70(21);
	sub_wire1(58, 22)    <= sub_wire70(22);
	sub_wire1(58, 23)    <= sub_wire70(23);
	sub_wire1(58, 24)    <= sub_wire70(24);
	sub_wire1(58, 25)    <= sub_wire70(25);
	sub_wire1(58, 26)    <= sub_wire70(26);
	sub_wire1(58, 27)    <= sub_wire70(27);
	sub_wire1(58, 28)    <= sub_wire70(28);
	sub_wire1(58, 29)    <= sub_wire70(29);
	sub_wire1(58, 30)    <= sub_wire70(30);
	sub_wire1(58, 31)    <= sub_wire70(31);
	sub_wire1(57, 0)    <= sub_wire71(0);
	sub_wire1(57, 1)    <= sub_wire71(1);
	sub_wire1(57, 2)    <= sub_wire71(2);
	sub_wire1(57, 3)    <= sub_wire71(3);
	sub_wire1(57, 4)    <= sub_wire71(4);
	sub_wire1(57, 5)    <= sub_wire71(5);
	sub_wire1(57, 6)    <= sub_wire71(6);
	sub_wire1(57, 7)    <= sub_wire71(7);
	sub_wire1(57, 8)    <= sub_wire71(8);
	sub_wire1(57, 9)    <= sub_wire71(9);
	sub_wire1(57, 10)    <= sub_wire71(10);
	sub_wire1(57, 11)    <= sub_wire71(11);
	sub_wire1(57, 12)    <= sub_wire71(12);
	sub_wire1(57, 13)    <= sub_wire71(13);
	sub_wire1(57, 14)    <= sub_wire71(14);
	sub_wire1(57, 15)    <= sub_wire71(15);
	sub_wire1(57, 16)    <= sub_wire71(16);
	sub_wire1(57, 17)    <= sub_wire71(17);
	sub_wire1(57, 18)    <= sub_wire71(18);
	sub_wire1(57, 19)    <= sub_wire71(19);
	sub_wire1(57, 20)    <= sub_wire71(20);
	sub_wire1(57, 21)    <= sub_wire71(21);
	sub_wire1(57, 22)    <= sub_wire71(22);
	sub_wire1(57, 23)    <= sub_wire71(23);
	sub_wire1(57, 24)    <= sub_wire71(24);
	sub_wire1(57, 25)    <= sub_wire71(25);
	sub_wire1(57, 26)    <= sub_wire71(26);
	sub_wire1(57, 27)    <= sub_wire71(27);
	sub_wire1(57, 28)    <= sub_wire71(28);
	sub_wire1(57, 29)    <= sub_wire71(29);
	sub_wire1(57, 30)    <= sub_wire71(30);
	sub_wire1(57, 31)    <= sub_wire71(31);
	sub_wire1(56, 0)    <= sub_wire72(0);
	sub_wire1(56, 1)    <= sub_wire72(1);
	sub_wire1(56, 2)    <= sub_wire72(2);
	sub_wire1(56, 3)    <= sub_wire72(3);
	sub_wire1(56, 4)    <= sub_wire72(4);
	sub_wire1(56, 5)    <= sub_wire72(5);
	sub_wire1(56, 6)    <= sub_wire72(6);
	sub_wire1(56, 7)    <= sub_wire72(7);
	sub_wire1(56, 8)    <= sub_wire72(8);
	sub_wire1(56, 9)    <= sub_wire72(9);
	sub_wire1(56, 10)    <= sub_wire72(10);
	sub_wire1(56, 11)    <= sub_wire72(11);
	sub_wire1(56, 12)    <= sub_wire72(12);
	sub_wire1(56, 13)    <= sub_wire72(13);
	sub_wire1(56, 14)    <= sub_wire72(14);
	sub_wire1(56, 15)    <= sub_wire72(15);
	sub_wire1(56, 16)    <= sub_wire72(16);
	sub_wire1(56, 17)    <= sub_wire72(17);
	sub_wire1(56, 18)    <= sub_wire72(18);
	sub_wire1(56, 19)    <= sub_wire72(19);
	sub_wire1(56, 20)    <= sub_wire72(20);
	sub_wire1(56, 21)    <= sub_wire72(21);
	sub_wire1(56, 22)    <= sub_wire72(22);
	sub_wire1(56, 23)    <= sub_wire72(23);
	sub_wire1(56, 24)    <= sub_wire72(24);
	sub_wire1(56, 25)    <= sub_wire72(25);
	sub_wire1(56, 26)    <= sub_wire72(26);
	sub_wire1(56, 27)    <= sub_wire72(27);
	sub_wire1(56, 28)    <= sub_wire72(28);
	sub_wire1(56, 29)    <= sub_wire72(29);
	sub_wire1(56, 30)    <= sub_wire72(30);
	sub_wire1(56, 31)    <= sub_wire72(31);
	sub_wire1(55, 0)    <= sub_wire73(0);
	sub_wire1(55, 1)    <= sub_wire73(1);
	sub_wire1(55, 2)    <= sub_wire73(2);
	sub_wire1(55, 3)    <= sub_wire73(3);
	sub_wire1(55, 4)    <= sub_wire73(4);
	sub_wire1(55, 5)    <= sub_wire73(5);
	sub_wire1(55, 6)    <= sub_wire73(6);
	sub_wire1(55, 7)    <= sub_wire73(7);
	sub_wire1(55, 8)    <= sub_wire73(8);
	sub_wire1(55, 9)    <= sub_wire73(9);
	sub_wire1(55, 10)    <= sub_wire73(10);
	sub_wire1(55, 11)    <= sub_wire73(11);
	sub_wire1(55, 12)    <= sub_wire73(12);
	sub_wire1(55, 13)    <= sub_wire73(13);
	sub_wire1(55, 14)    <= sub_wire73(14);
	sub_wire1(55, 15)    <= sub_wire73(15);
	sub_wire1(55, 16)    <= sub_wire73(16);
	sub_wire1(55, 17)    <= sub_wire73(17);
	sub_wire1(55, 18)    <= sub_wire73(18);
	sub_wire1(55, 19)    <= sub_wire73(19);
	sub_wire1(55, 20)    <= sub_wire73(20);
	sub_wire1(55, 21)    <= sub_wire73(21);
	sub_wire1(55, 22)    <= sub_wire73(22);
	sub_wire1(55, 23)    <= sub_wire73(23);
	sub_wire1(55, 24)    <= sub_wire73(24);
	sub_wire1(55, 25)    <= sub_wire73(25);
	sub_wire1(55, 26)    <= sub_wire73(26);
	sub_wire1(55, 27)    <= sub_wire73(27);
	sub_wire1(55, 28)    <= sub_wire73(28);
	sub_wire1(55, 29)    <= sub_wire73(29);
	sub_wire1(55, 30)    <= sub_wire73(30);
	sub_wire1(55, 31)    <= sub_wire73(31);
	sub_wire1(54, 0)    <= sub_wire74(0);
	sub_wire1(54, 1)    <= sub_wire74(1);
	sub_wire1(54, 2)    <= sub_wire74(2);
	sub_wire1(54, 3)    <= sub_wire74(3);
	sub_wire1(54, 4)    <= sub_wire74(4);
	sub_wire1(54, 5)    <= sub_wire74(5);
	sub_wire1(54, 6)    <= sub_wire74(6);
	sub_wire1(54, 7)    <= sub_wire74(7);
	sub_wire1(54, 8)    <= sub_wire74(8);
	sub_wire1(54, 9)    <= sub_wire74(9);
	sub_wire1(54, 10)    <= sub_wire74(10);
	sub_wire1(54, 11)    <= sub_wire74(11);
	sub_wire1(54, 12)    <= sub_wire74(12);
	sub_wire1(54, 13)    <= sub_wire74(13);
	sub_wire1(54, 14)    <= sub_wire74(14);
	sub_wire1(54, 15)    <= sub_wire74(15);
	sub_wire1(54, 16)    <= sub_wire74(16);
	sub_wire1(54, 17)    <= sub_wire74(17);
	sub_wire1(54, 18)    <= sub_wire74(18);
	sub_wire1(54, 19)    <= sub_wire74(19);
	sub_wire1(54, 20)    <= sub_wire74(20);
	sub_wire1(54, 21)    <= sub_wire74(21);
	sub_wire1(54, 22)    <= sub_wire74(22);
	sub_wire1(54, 23)    <= sub_wire74(23);
	sub_wire1(54, 24)    <= sub_wire74(24);
	sub_wire1(54, 25)    <= sub_wire74(25);
	sub_wire1(54, 26)    <= sub_wire74(26);
	sub_wire1(54, 27)    <= sub_wire74(27);
	sub_wire1(54, 28)    <= sub_wire74(28);
	sub_wire1(54, 29)    <= sub_wire74(29);
	sub_wire1(54, 30)    <= sub_wire74(30);
	sub_wire1(54, 31)    <= sub_wire74(31);
	sub_wire1(53, 0)    <= sub_wire75(0);
	sub_wire1(53, 1)    <= sub_wire75(1);
	sub_wire1(53, 2)    <= sub_wire75(2);
	sub_wire1(53, 3)    <= sub_wire75(3);
	sub_wire1(53, 4)    <= sub_wire75(4);
	sub_wire1(53, 5)    <= sub_wire75(5);
	sub_wire1(53, 6)    <= sub_wire75(6);
	sub_wire1(53, 7)    <= sub_wire75(7);
	sub_wire1(53, 8)    <= sub_wire75(8);
	sub_wire1(53, 9)    <= sub_wire75(9);
	sub_wire1(53, 10)    <= sub_wire75(10);
	sub_wire1(53, 11)    <= sub_wire75(11);
	sub_wire1(53, 12)    <= sub_wire75(12);
	sub_wire1(53, 13)    <= sub_wire75(13);
	sub_wire1(53, 14)    <= sub_wire75(14);
	sub_wire1(53, 15)    <= sub_wire75(15);
	sub_wire1(53, 16)    <= sub_wire75(16);
	sub_wire1(53, 17)    <= sub_wire75(17);
	sub_wire1(53, 18)    <= sub_wire75(18);
	sub_wire1(53, 19)    <= sub_wire75(19);
	sub_wire1(53, 20)    <= sub_wire75(20);
	sub_wire1(53, 21)    <= sub_wire75(21);
	sub_wire1(53, 22)    <= sub_wire75(22);
	sub_wire1(53, 23)    <= sub_wire75(23);
	sub_wire1(53, 24)    <= sub_wire75(24);
	sub_wire1(53, 25)    <= sub_wire75(25);
	sub_wire1(53, 26)    <= sub_wire75(26);
	sub_wire1(53, 27)    <= sub_wire75(27);
	sub_wire1(53, 28)    <= sub_wire75(28);
	sub_wire1(53, 29)    <= sub_wire75(29);
	sub_wire1(53, 30)    <= sub_wire75(30);
	sub_wire1(53, 31)    <= sub_wire75(31);
	sub_wire1(52, 0)    <= sub_wire76(0);
	sub_wire1(52, 1)    <= sub_wire76(1);
	sub_wire1(52, 2)    <= sub_wire76(2);
	sub_wire1(52, 3)    <= sub_wire76(3);
	sub_wire1(52, 4)    <= sub_wire76(4);
	sub_wire1(52, 5)    <= sub_wire76(5);
	sub_wire1(52, 6)    <= sub_wire76(6);
	sub_wire1(52, 7)    <= sub_wire76(7);
	sub_wire1(52, 8)    <= sub_wire76(8);
	sub_wire1(52, 9)    <= sub_wire76(9);
	sub_wire1(52, 10)    <= sub_wire76(10);
	sub_wire1(52, 11)    <= sub_wire76(11);
	sub_wire1(52, 12)    <= sub_wire76(12);
	sub_wire1(52, 13)    <= sub_wire76(13);
	sub_wire1(52, 14)    <= sub_wire76(14);
	sub_wire1(52, 15)    <= sub_wire76(15);
	sub_wire1(52, 16)    <= sub_wire76(16);
	sub_wire1(52, 17)    <= sub_wire76(17);
	sub_wire1(52, 18)    <= sub_wire76(18);
	sub_wire1(52, 19)    <= sub_wire76(19);
	sub_wire1(52, 20)    <= sub_wire76(20);
	sub_wire1(52, 21)    <= sub_wire76(21);
	sub_wire1(52, 22)    <= sub_wire76(22);
	sub_wire1(52, 23)    <= sub_wire76(23);
	sub_wire1(52, 24)    <= sub_wire76(24);
	sub_wire1(52, 25)    <= sub_wire76(25);
	sub_wire1(52, 26)    <= sub_wire76(26);
	sub_wire1(52, 27)    <= sub_wire76(27);
	sub_wire1(52, 28)    <= sub_wire76(28);
	sub_wire1(52, 29)    <= sub_wire76(29);
	sub_wire1(52, 30)    <= sub_wire76(30);
	sub_wire1(52, 31)    <= sub_wire76(31);
	sub_wire1(51, 0)    <= sub_wire77(0);
	sub_wire1(51, 1)    <= sub_wire77(1);
	sub_wire1(51, 2)    <= sub_wire77(2);
	sub_wire1(51, 3)    <= sub_wire77(3);
	sub_wire1(51, 4)    <= sub_wire77(4);
	sub_wire1(51, 5)    <= sub_wire77(5);
	sub_wire1(51, 6)    <= sub_wire77(6);
	sub_wire1(51, 7)    <= sub_wire77(7);
	sub_wire1(51, 8)    <= sub_wire77(8);
	sub_wire1(51, 9)    <= sub_wire77(9);
	sub_wire1(51, 10)    <= sub_wire77(10);
	sub_wire1(51, 11)    <= sub_wire77(11);
	sub_wire1(51, 12)    <= sub_wire77(12);
	sub_wire1(51, 13)    <= sub_wire77(13);
	sub_wire1(51, 14)    <= sub_wire77(14);
	sub_wire1(51, 15)    <= sub_wire77(15);
	sub_wire1(51, 16)    <= sub_wire77(16);
	sub_wire1(51, 17)    <= sub_wire77(17);
	sub_wire1(51, 18)    <= sub_wire77(18);
	sub_wire1(51, 19)    <= sub_wire77(19);
	sub_wire1(51, 20)    <= sub_wire77(20);
	sub_wire1(51, 21)    <= sub_wire77(21);
	sub_wire1(51, 22)    <= sub_wire77(22);
	sub_wire1(51, 23)    <= sub_wire77(23);
	sub_wire1(51, 24)    <= sub_wire77(24);
	sub_wire1(51, 25)    <= sub_wire77(25);
	sub_wire1(51, 26)    <= sub_wire77(26);
	sub_wire1(51, 27)    <= sub_wire77(27);
	sub_wire1(51, 28)    <= sub_wire77(28);
	sub_wire1(51, 29)    <= sub_wire77(29);
	sub_wire1(51, 30)    <= sub_wire77(30);
	sub_wire1(51, 31)    <= sub_wire77(31);
	sub_wire1(50, 0)    <= sub_wire78(0);
	sub_wire1(50, 1)    <= sub_wire78(1);
	sub_wire1(50, 2)    <= sub_wire78(2);
	sub_wire1(50, 3)    <= sub_wire78(3);
	sub_wire1(50, 4)    <= sub_wire78(4);
	sub_wire1(50, 5)    <= sub_wire78(5);
	sub_wire1(50, 6)    <= sub_wire78(6);
	sub_wire1(50, 7)    <= sub_wire78(7);
	sub_wire1(50, 8)    <= sub_wire78(8);
	sub_wire1(50, 9)    <= sub_wire78(9);
	sub_wire1(50, 10)    <= sub_wire78(10);
	sub_wire1(50, 11)    <= sub_wire78(11);
	sub_wire1(50, 12)    <= sub_wire78(12);
	sub_wire1(50, 13)    <= sub_wire78(13);
	sub_wire1(50, 14)    <= sub_wire78(14);
	sub_wire1(50, 15)    <= sub_wire78(15);
	sub_wire1(50, 16)    <= sub_wire78(16);
	sub_wire1(50, 17)    <= sub_wire78(17);
	sub_wire1(50, 18)    <= sub_wire78(18);
	sub_wire1(50, 19)    <= sub_wire78(19);
	sub_wire1(50, 20)    <= sub_wire78(20);
	sub_wire1(50, 21)    <= sub_wire78(21);
	sub_wire1(50, 22)    <= sub_wire78(22);
	sub_wire1(50, 23)    <= sub_wire78(23);
	sub_wire1(50, 24)    <= sub_wire78(24);
	sub_wire1(50, 25)    <= sub_wire78(25);
	sub_wire1(50, 26)    <= sub_wire78(26);
	sub_wire1(50, 27)    <= sub_wire78(27);
	sub_wire1(50, 28)    <= sub_wire78(28);
	sub_wire1(50, 29)    <= sub_wire78(29);
	sub_wire1(50, 30)    <= sub_wire78(30);
	sub_wire1(50, 31)    <= sub_wire78(31);
	sub_wire1(49, 0)    <= sub_wire79(0);
	sub_wire1(49, 1)    <= sub_wire79(1);
	sub_wire1(49, 2)    <= sub_wire79(2);
	sub_wire1(49, 3)    <= sub_wire79(3);
	sub_wire1(49, 4)    <= sub_wire79(4);
	sub_wire1(49, 5)    <= sub_wire79(5);
	sub_wire1(49, 6)    <= sub_wire79(6);
	sub_wire1(49, 7)    <= sub_wire79(7);
	sub_wire1(49, 8)    <= sub_wire79(8);
	sub_wire1(49, 9)    <= sub_wire79(9);
	sub_wire1(49, 10)    <= sub_wire79(10);
	sub_wire1(49, 11)    <= sub_wire79(11);
	sub_wire1(49, 12)    <= sub_wire79(12);
	sub_wire1(49, 13)    <= sub_wire79(13);
	sub_wire1(49, 14)    <= sub_wire79(14);
	sub_wire1(49, 15)    <= sub_wire79(15);
	sub_wire1(49, 16)    <= sub_wire79(16);
	sub_wire1(49, 17)    <= sub_wire79(17);
	sub_wire1(49, 18)    <= sub_wire79(18);
	sub_wire1(49, 19)    <= sub_wire79(19);
	sub_wire1(49, 20)    <= sub_wire79(20);
	sub_wire1(49, 21)    <= sub_wire79(21);
	sub_wire1(49, 22)    <= sub_wire79(22);
	sub_wire1(49, 23)    <= sub_wire79(23);
	sub_wire1(49, 24)    <= sub_wire79(24);
	sub_wire1(49, 25)    <= sub_wire79(25);
	sub_wire1(49, 26)    <= sub_wire79(26);
	sub_wire1(49, 27)    <= sub_wire79(27);
	sub_wire1(49, 28)    <= sub_wire79(28);
	sub_wire1(49, 29)    <= sub_wire79(29);
	sub_wire1(49, 30)    <= sub_wire79(30);
	sub_wire1(49, 31)    <= sub_wire79(31);
	sub_wire1(48, 0)    <= sub_wire80(0);
	sub_wire1(48, 1)    <= sub_wire80(1);
	sub_wire1(48, 2)    <= sub_wire80(2);
	sub_wire1(48, 3)    <= sub_wire80(3);
	sub_wire1(48, 4)    <= sub_wire80(4);
	sub_wire1(48, 5)    <= sub_wire80(5);
	sub_wire1(48, 6)    <= sub_wire80(6);
	sub_wire1(48, 7)    <= sub_wire80(7);
	sub_wire1(48, 8)    <= sub_wire80(8);
	sub_wire1(48, 9)    <= sub_wire80(9);
	sub_wire1(48, 10)    <= sub_wire80(10);
	sub_wire1(48, 11)    <= sub_wire80(11);
	sub_wire1(48, 12)    <= sub_wire80(12);
	sub_wire1(48, 13)    <= sub_wire80(13);
	sub_wire1(48, 14)    <= sub_wire80(14);
	sub_wire1(48, 15)    <= sub_wire80(15);
	sub_wire1(48, 16)    <= sub_wire80(16);
	sub_wire1(48, 17)    <= sub_wire80(17);
	sub_wire1(48, 18)    <= sub_wire80(18);
	sub_wire1(48, 19)    <= sub_wire80(19);
	sub_wire1(48, 20)    <= sub_wire80(20);
	sub_wire1(48, 21)    <= sub_wire80(21);
	sub_wire1(48, 22)    <= sub_wire80(22);
	sub_wire1(48, 23)    <= sub_wire80(23);
	sub_wire1(48, 24)    <= sub_wire80(24);
	sub_wire1(48, 25)    <= sub_wire80(25);
	sub_wire1(48, 26)    <= sub_wire80(26);
	sub_wire1(48, 27)    <= sub_wire80(27);
	sub_wire1(48, 28)    <= sub_wire80(28);
	sub_wire1(48, 29)    <= sub_wire80(29);
	sub_wire1(48, 30)    <= sub_wire80(30);
	sub_wire1(48, 31)    <= sub_wire80(31);
	sub_wire1(47, 0)    <= sub_wire81(0);
	sub_wire1(47, 1)    <= sub_wire81(1);
	sub_wire1(47, 2)    <= sub_wire81(2);
	sub_wire1(47, 3)    <= sub_wire81(3);
	sub_wire1(47, 4)    <= sub_wire81(4);
	sub_wire1(47, 5)    <= sub_wire81(5);
	sub_wire1(47, 6)    <= sub_wire81(6);
	sub_wire1(47, 7)    <= sub_wire81(7);
	sub_wire1(47, 8)    <= sub_wire81(8);
	sub_wire1(47, 9)    <= sub_wire81(9);
	sub_wire1(47, 10)    <= sub_wire81(10);
	sub_wire1(47, 11)    <= sub_wire81(11);
	sub_wire1(47, 12)    <= sub_wire81(12);
	sub_wire1(47, 13)    <= sub_wire81(13);
	sub_wire1(47, 14)    <= sub_wire81(14);
	sub_wire1(47, 15)    <= sub_wire81(15);
	sub_wire1(47, 16)    <= sub_wire81(16);
	sub_wire1(47, 17)    <= sub_wire81(17);
	sub_wire1(47, 18)    <= sub_wire81(18);
	sub_wire1(47, 19)    <= sub_wire81(19);
	sub_wire1(47, 20)    <= sub_wire81(20);
	sub_wire1(47, 21)    <= sub_wire81(21);
	sub_wire1(47, 22)    <= sub_wire81(22);
	sub_wire1(47, 23)    <= sub_wire81(23);
	sub_wire1(47, 24)    <= sub_wire81(24);
	sub_wire1(47, 25)    <= sub_wire81(25);
	sub_wire1(47, 26)    <= sub_wire81(26);
	sub_wire1(47, 27)    <= sub_wire81(27);
	sub_wire1(47, 28)    <= sub_wire81(28);
	sub_wire1(47, 29)    <= sub_wire81(29);
	sub_wire1(47, 30)    <= sub_wire81(30);
	sub_wire1(47, 31)    <= sub_wire81(31);
	sub_wire1(46, 0)    <= sub_wire82(0);
	sub_wire1(46, 1)    <= sub_wire82(1);
	sub_wire1(46, 2)    <= sub_wire82(2);
	sub_wire1(46, 3)    <= sub_wire82(3);
	sub_wire1(46, 4)    <= sub_wire82(4);
	sub_wire1(46, 5)    <= sub_wire82(5);
	sub_wire1(46, 6)    <= sub_wire82(6);
	sub_wire1(46, 7)    <= sub_wire82(7);
	sub_wire1(46, 8)    <= sub_wire82(8);
	sub_wire1(46, 9)    <= sub_wire82(9);
	sub_wire1(46, 10)    <= sub_wire82(10);
	sub_wire1(46, 11)    <= sub_wire82(11);
	sub_wire1(46, 12)    <= sub_wire82(12);
	sub_wire1(46, 13)    <= sub_wire82(13);
	sub_wire1(46, 14)    <= sub_wire82(14);
	sub_wire1(46, 15)    <= sub_wire82(15);
	sub_wire1(46, 16)    <= sub_wire82(16);
	sub_wire1(46, 17)    <= sub_wire82(17);
	sub_wire1(46, 18)    <= sub_wire82(18);
	sub_wire1(46, 19)    <= sub_wire82(19);
	sub_wire1(46, 20)    <= sub_wire82(20);
	sub_wire1(46, 21)    <= sub_wire82(21);
	sub_wire1(46, 22)    <= sub_wire82(22);
	sub_wire1(46, 23)    <= sub_wire82(23);
	sub_wire1(46, 24)    <= sub_wire82(24);
	sub_wire1(46, 25)    <= sub_wire82(25);
	sub_wire1(46, 26)    <= sub_wire82(26);
	sub_wire1(46, 27)    <= sub_wire82(27);
	sub_wire1(46, 28)    <= sub_wire82(28);
	sub_wire1(46, 29)    <= sub_wire82(29);
	sub_wire1(46, 30)    <= sub_wire82(30);
	sub_wire1(46, 31)    <= sub_wire82(31);
	sub_wire1(45, 0)    <= sub_wire83(0);
	sub_wire1(45, 1)    <= sub_wire83(1);
	sub_wire1(45, 2)    <= sub_wire83(2);
	sub_wire1(45, 3)    <= sub_wire83(3);
	sub_wire1(45, 4)    <= sub_wire83(4);
	sub_wire1(45, 5)    <= sub_wire83(5);
	sub_wire1(45, 6)    <= sub_wire83(6);
	sub_wire1(45, 7)    <= sub_wire83(7);
	sub_wire1(45, 8)    <= sub_wire83(8);
	sub_wire1(45, 9)    <= sub_wire83(9);
	sub_wire1(45, 10)    <= sub_wire83(10);
	sub_wire1(45, 11)    <= sub_wire83(11);
	sub_wire1(45, 12)    <= sub_wire83(12);
	sub_wire1(45, 13)    <= sub_wire83(13);
	sub_wire1(45, 14)    <= sub_wire83(14);
	sub_wire1(45, 15)    <= sub_wire83(15);
	sub_wire1(45, 16)    <= sub_wire83(16);
	sub_wire1(45, 17)    <= sub_wire83(17);
	sub_wire1(45, 18)    <= sub_wire83(18);
	sub_wire1(45, 19)    <= sub_wire83(19);
	sub_wire1(45, 20)    <= sub_wire83(20);
	sub_wire1(45, 21)    <= sub_wire83(21);
	sub_wire1(45, 22)    <= sub_wire83(22);
	sub_wire1(45, 23)    <= sub_wire83(23);
	sub_wire1(45, 24)    <= sub_wire83(24);
	sub_wire1(45, 25)    <= sub_wire83(25);
	sub_wire1(45, 26)    <= sub_wire83(26);
	sub_wire1(45, 27)    <= sub_wire83(27);
	sub_wire1(45, 28)    <= sub_wire83(28);
	sub_wire1(45, 29)    <= sub_wire83(29);
	sub_wire1(45, 30)    <= sub_wire83(30);
	sub_wire1(45, 31)    <= sub_wire83(31);
	sub_wire1(44, 0)    <= sub_wire84(0);
	sub_wire1(44, 1)    <= sub_wire84(1);
	sub_wire1(44, 2)    <= sub_wire84(2);
	sub_wire1(44, 3)    <= sub_wire84(3);
	sub_wire1(44, 4)    <= sub_wire84(4);
	sub_wire1(44, 5)    <= sub_wire84(5);
	sub_wire1(44, 6)    <= sub_wire84(6);
	sub_wire1(44, 7)    <= sub_wire84(7);
	sub_wire1(44, 8)    <= sub_wire84(8);
	sub_wire1(44, 9)    <= sub_wire84(9);
	sub_wire1(44, 10)    <= sub_wire84(10);
	sub_wire1(44, 11)    <= sub_wire84(11);
	sub_wire1(44, 12)    <= sub_wire84(12);
	sub_wire1(44, 13)    <= sub_wire84(13);
	sub_wire1(44, 14)    <= sub_wire84(14);
	sub_wire1(44, 15)    <= sub_wire84(15);
	sub_wire1(44, 16)    <= sub_wire84(16);
	sub_wire1(44, 17)    <= sub_wire84(17);
	sub_wire1(44, 18)    <= sub_wire84(18);
	sub_wire1(44, 19)    <= sub_wire84(19);
	sub_wire1(44, 20)    <= sub_wire84(20);
	sub_wire1(44, 21)    <= sub_wire84(21);
	sub_wire1(44, 22)    <= sub_wire84(22);
	sub_wire1(44, 23)    <= sub_wire84(23);
	sub_wire1(44, 24)    <= sub_wire84(24);
	sub_wire1(44, 25)    <= sub_wire84(25);
	sub_wire1(44, 26)    <= sub_wire84(26);
	sub_wire1(44, 27)    <= sub_wire84(27);
	sub_wire1(44, 28)    <= sub_wire84(28);
	sub_wire1(44, 29)    <= sub_wire84(29);
	sub_wire1(44, 30)    <= sub_wire84(30);
	sub_wire1(44, 31)    <= sub_wire84(31);
	sub_wire1(43, 0)    <= sub_wire85(0);
	sub_wire1(43, 1)    <= sub_wire85(1);
	sub_wire1(43, 2)    <= sub_wire85(2);
	sub_wire1(43, 3)    <= sub_wire85(3);
	sub_wire1(43, 4)    <= sub_wire85(4);
	sub_wire1(43, 5)    <= sub_wire85(5);
	sub_wire1(43, 6)    <= sub_wire85(6);
	sub_wire1(43, 7)    <= sub_wire85(7);
	sub_wire1(43, 8)    <= sub_wire85(8);
	sub_wire1(43, 9)    <= sub_wire85(9);
	sub_wire1(43, 10)    <= sub_wire85(10);
	sub_wire1(43, 11)    <= sub_wire85(11);
	sub_wire1(43, 12)    <= sub_wire85(12);
	sub_wire1(43, 13)    <= sub_wire85(13);
	sub_wire1(43, 14)    <= sub_wire85(14);
	sub_wire1(43, 15)    <= sub_wire85(15);
	sub_wire1(43, 16)    <= sub_wire85(16);
	sub_wire1(43, 17)    <= sub_wire85(17);
	sub_wire1(43, 18)    <= sub_wire85(18);
	sub_wire1(43, 19)    <= sub_wire85(19);
	sub_wire1(43, 20)    <= sub_wire85(20);
	sub_wire1(43, 21)    <= sub_wire85(21);
	sub_wire1(43, 22)    <= sub_wire85(22);
	sub_wire1(43, 23)    <= sub_wire85(23);
	sub_wire1(43, 24)    <= sub_wire85(24);
	sub_wire1(43, 25)    <= sub_wire85(25);
	sub_wire1(43, 26)    <= sub_wire85(26);
	sub_wire1(43, 27)    <= sub_wire85(27);
	sub_wire1(43, 28)    <= sub_wire85(28);
	sub_wire1(43, 29)    <= sub_wire85(29);
	sub_wire1(43, 30)    <= sub_wire85(30);
	sub_wire1(43, 31)    <= sub_wire85(31);
	sub_wire1(42, 0)    <= sub_wire86(0);
	sub_wire1(42, 1)    <= sub_wire86(1);
	sub_wire1(42, 2)    <= sub_wire86(2);
	sub_wire1(42, 3)    <= sub_wire86(3);
	sub_wire1(42, 4)    <= sub_wire86(4);
	sub_wire1(42, 5)    <= sub_wire86(5);
	sub_wire1(42, 6)    <= sub_wire86(6);
	sub_wire1(42, 7)    <= sub_wire86(7);
	sub_wire1(42, 8)    <= sub_wire86(8);
	sub_wire1(42, 9)    <= sub_wire86(9);
	sub_wire1(42, 10)    <= sub_wire86(10);
	sub_wire1(42, 11)    <= sub_wire86(11);
	sub_wire1(42, 12)    <= sub_wire86(12);
	sub_wire1(42, 13)    <= sub_wire86(13);
	sub_wire1(42, 14)    <= sub_wire86(14);
	sub_wire1(42, 15)    <= sub_wire86(15);
	sub_wire1(42, 16)    <= sub_wire86(16);
	sub_wire1(42, 17)    <= sub_wire86(17);
	sub_wire1(42, 18)    <= sub_wire86(18);
	sub_wire1(42, 19)    <= sub_wire86(19);
	sub_wire1(42, 20)    <= sub_wire86(20);
	sub_wire1(42, 21)    <= sub_wire86(21);
	sub_wire1(42, 22)    <= sub_wire86(22);
	sub_wire1(42, 23)    <= sub_wire86(23);
	sub_wire1(42, 24)    <= sub_wire86(24);
	sub_wire1(42, 25)    <= sub_wire86(25);
	sub_wire1(42, 26)    <= sub_wire86(26);
	sub_wire1(42, 27)    <= sub_wire86(27);
	sub_wire1(42, 28)    <= sub_wire86(28);
	sub_wire1(42, 29)    <= sub_wire86(29);
	sub_wire1(42, 30)    <= sub_wire86(30);
	sub_wire1(42, 31)    <= sub_wire86(31);
	sub_wire1(41, 0)    <= sub_wire87(0);
	sub_wire1(41, 1)    <= sub_wire87(1);
	sub_wire1(41, 2)    <= sub_wire87(2);
	sub_wire1(41, 3)    <= sub_wire87(3);
	sub_wire1(41, 4)    <= sub_wire87(4);
	sub_wire1(41, 5)    <= sub_wire87(5);
	sub_wire1(41, 6)    <= sub_wire87(6);
	sub_wire1(41, 7)    <= sub_wire87(7);
	sub_wire1(41, 8)    <= sub_wire87(8);
	sub_wire1(41, 9)    <= sub_wire87(9);
	sub_wire1(41, 10)    <= sub_wire87(10);
	sub_wire1(41, 11)    <= sub_wire87(11);
	sub_wire1(41, 12)    <= sub_wire87(12);
	sub_wire1(41, 13)    <= sub_wire87(13);
	sub_wire1(41, 14)    <= sub_wire87(14);
	sub_wire1(41, 15)    <= sub_wire87(15);
	sub_wire1(41, 16)    <= sub_wire87(16);
	sub_wire1(41, 17)    <= sub_wire87(17);
	sub_wire1(41, 18)    <= sub_wire87(18);
	sub_wire1(41, 19)    <= sub_wire87(19);
	sub_wire1(41, 20)    <= sub_wire87(20);
	sub_wire1(41, 21)    <= sub_wire87(21);
	sub_wire1(41, 22)    <= sub_wire87(22);
	sub_wire1(41, 23)    <= sub_wire87(23);
	sub_wire1(41, 24)    <= sub_wire87(24);
	sub_wire1(41, 25)    <= sub_wire87(25);
	sub_wire1(41, 26)    <= sub_wire87(26);
	sub_wire1(41, 27)    <= sub_wire87(27);
	sub_wire1(41, 28)    <= sub_wire87(28);
	sub_wire1(41, 29)    <= sub_wire87(29);
	sub_wire1(41, 30)    <= sub_wire87(30);
	sub_wire1(41, 31)    <= sub_wire87(31);
	sub_wire1(40, 0)    <= sub_wire88(0);
	sub_wire1(40, 1)    <= sub_wire88(1);
	sub_wire1(40, 2)    <= sub_wire88(2);
	sub_wire1(40, 3)    <= sub_wire88(3);
	sub_wire1(40, 4)    <= sub_wire88(4);
	sub_wire1(40, 5)    <= sub_wire88(5);
	sub_wire1(40, 6)    <= sub_wire88(6);
	sub_wire1(40, 7)    <= sub_wire88(7);
	sub_wire1(40, 8)    <= sub_wire88(8);
	sub_wire1(40, 9)    <= sub_wire88(9);
	sub_wire1(40, 10)    <= sub_wire88(10);
	sub_wire1(40, 11)    <= sub_wire88(11);
	sub_wire1(40, 12)    <= sub_wire88(12);
	sub_wire1(40, 13)    <= sub_wire88(13);
	sub_wire1(40, 14)    <= sub_wire88(14);
	sub_wire1(40, 15)    <= sub_wire88(15);
	sub_wire1(40, 16)    <= sub_wire88(16);
	sub_wire1(40, 17)    <= sub_wire88(17);
	sub_wire1(40, 18)    <= sub_wire88(18);
	sub_wire1(40, 19)    <= sub_wire88(19);
	sub_wire1(40, 20)    <= sub_wire88(20);
	sub_wire1(40, 21)    <= sub_wire88(21);
	sub_wire1(40, 22)    <= sub_wire88(22);
	sub_wire1(40, 23)    <= sub_wire88(23);
	sub_wire1(40, 24)    <= sub_wire88(24);
	sub_wire1(40, 25)    <= sub_wire88(25);
	sub_wire1(40, 26)    <= sub_wire88(26);
	sub_wire1(40, 27)    <= sub_wire88(27);
	sub_wire1(40, 28)    <= sub_wire88(28);
	sub_wire1(40, 29)    <= sub_wire88(29);
	sub_wire1(40, 30)    <= sub_wire88(30);
	sub_wire1(40, 31)    <= sub_wire88(31);
	sub_wire1(39, 0)    <= sub_wire89(0);
	sub_wire1(39, 1)    <= sub_wire89(1);
	sub_wire1(39, 2)    <= sub_wire89(2);
	sub_wire1(39, 3)    <= sub_wire89(3);
	sub_wire1(39, 4)    <= sub_wire89(4);
	sub_wire1(39, 5)    <= sub_wire89(5);
	sub_wire1(39, 6)    <= sub_wire89(6);
	sub_wire1(39, 7)    <= sub_wire89(7);
	sub_wire1(39, 8)    <= sub_wire89(8);
	sub_wire1(39, 9)    <= sub_wire89(9);
	sub_wire1(39, 10)    <= sub_wire89(10);
	sub_wire1(39, 11)    <= sub_wire89(11);
	sub_wire1(39, 12)    <= sub_wire89(12);
	sub_wire1(39, 13)    <= sub_wire89(13);
	sub_wire1(39, 14)    <= sub_wire89(14);
	sub_wire1(39, 15)    <= sub_wire89(15);
	sub_wire1(39, 16)    <= sub_wire89(16);
	sub_wire1(39, 17)    <= sub_wire89(17);
	sub_wire1(39, 18)    <= sub_wire89(18);
	sub_wire1(39, 19)    <= sub_wire89(19);
	sub_wire1(39, 20)    <= sub_wire89(20);
	sub_wire1(39, 21)    <= sub_wire89(21);
	sub_wire1(39, 22)    <= sub_wire89(22);
	sub_wire1(39, 23)    <= sub_wire89(23);
	sub_wire1(39, 24)    <= sub_wire89(24);
	sub_wire1(39, 25)    <= sub_wire89(25);
	sub_wire1(39, 26)    <= sub_wire89(26);
	sub_wire1(39, 27)    <= sub_wire89(27);
	sub_wire1(39, 28)    <= sub_wire89(28);
	sub_wire1(39, 29)    <= sub_wire89(29);
	sub_wire1(39, 30)    <= sub_wire89(30);
	sub_wire1(39, 31)    <= sub_wire89(31);
	sub_wire1(38, 0)    <= sub_wire90(0);
	sub_wire1(38, 1)    <= sub_wire90(1);
	sub_wire1(38, 2)    <= sub_wire90(2);
	sub_wire1(38, 3)    <= sub_wire90(3);
	sub_wire1(38, 4)    <= sub_wire90(4);
	sub_wire1(38, 5)    <= sub_wire90(5);
	sub_wire1(38, 6)    <= sub_wire90(6);
	sub_wire1(38, 7)    <= sub_wire90(7);
	sub_wire1(38, 8)    <= sub_wire90(8);
	sub_wire1(38, 9)    <= sub_wire90(9);
	sub_wire1(38, 10)    <= sub_wire90(10);
	sub_wire1(38, 11)    <= sub_wire90(11);
	sub_wire1(38, 12)    <= sub_wire90(12);
	sub_wire1(38, 13)    <= sub_wire90(13);
	sub_wire1(38, 14)    <= sub_wire90(14);
	sub_wire1(38, 15)    <= sub_wire90(15);
	sub_wire1(38, 16)    <= sub_wire90(16);
	sub_wire1(38, 17)    <= sub_wire90(17);
	sub_wire1(38, 18)    <= sub_wire90(18);
	sub_wire1(38, 19)    <= sub_wire90(19);
	sub_wire1(38, 20)    <= sub_wire90(20);
	sub_wire1(38, 21)    <= sub_wire90(21);
	sub_wire1(38, 22)    <= sub_wire90(22);
	sub_wire1(38, 23)    <= sub_wire90(23);
	sub_wire1(38, 24)    <= sub_wire90(24);
	sub_wire1(38, 25)    <= sub_wire90(25);
	sub_wire1(38, 26)    <= sub_wire90(26);
	sub_wire1(38, 27)    <= sub_wire90(27);
	sub_wire1(38, 28)    <= sub_wire90(28);
	sub_wire1(38, 29)    <= sub_wire90(29);
	sub_wire1(38, 30)    <= sub_wire90(30);
	sub_wire1(38, 31)    <= sub_wire90(31);
	sub_wire1(37, 0)    <= sub_wire91(0);
	sub_wire1(37, 1)    <= sub_wire91(1);
	sub_wire1(37, 2)    <= sub_wire91(2);
	sub_wire1(37, 3)    <= sub_wire91(3);
	sub_wire1(37, 4)    <= sub_wire91(4);
	sub_wire1(37, 5)    <= sub_wire91(5);
	sub_wire1(37, 6)    <= sub_wire91(6);
	sub_wire1(37, 7)    <= sub_wire91(7);
	sub_wire1(37, 8)    <= sub_wire91(8);
	sub_wire1(37, 9)    <= sub_wire91(9);
	sub_wire1(37, 10)    <= sub_wire91(10);
	sub_wire1(37, 11)    <= sub_wire91(11);
	sub_wire1(37, 12)    <= sub_wire91(12);
	sub_wire1(37, 13)    <= sub_wire91(13);
	sub_wire1(37, 14)    <= sub_wire91(14);
	sub_wire1(37, 15)    <= sub_wire91(15);
	sub_wire1(37, 16)    <= sub_wire91(16);
	sub_wire1(37, 17)    <= sub_wire91(17);
	sub_wire1(37, 18)    <= sub_wire91(18);
	sub_wire1(37, 19)    <= sub_wire91(19);
	sub_wire1(37, 20)    <= sub_wire91(20);
	sub_wire1(37, 21)    <= sub_wire91(21);
	sub_wire1(37, 22)    <= sub_wire91(22);
	sub_wire1(37, 23)    <= sub_wire91(23);
	sub_wire1(37, 24)    <= sub_wire91(24);
	sub_wire1(37, 25)    <= sub_wire91(25);
	sub_wire1(37, 26)    <= sub_wire91(26);
	sub_wire1(37, 27)    <= sub_wire91(27);
	sub_wire1(37, 28)    <= sub_wire91(28);
	sub_wire1(37, 29)    <= sub_wire91(29);
	sub_wire1(37, 30)    <= sub_wire91(30);
	sub_wire1(37, 31)    <= sub_wire91(31);
	sub_wire1(36, 0)    <= sub_wire92(0);
	sub_wire1(36, 1)    <= sub_wire92(1);
	sub_wire1(36, 2)    <= sub_wire92(2);
	sub_wire1(36, 3)    <= sub_wire92(3);
	sub_wire1(36, 4)    <= sub_wire92(4);
	sub_wire1(36, 5)    <= sub_wire92(5);
	sub_wire1(36, 6)    <= sub_wire92(6);
	sub_wire1(36, 7)    <= sub_wire92(7);
	sub_wire1(36, 8)    <= sub_wire92(8);
	sub_wire1(36, 9)    <= sub_wire92(9);
	sub_wire1(36, 10)    <= sub_wire92(10);
	sub_wire1(36, 11)    <= sub_wire92(11);
	sub_wire1(36, 12)    <= sub_wire92(12);
	sub_wire1(36, 13)    <= sub_wire92(13);
	sub_wire1(36, 14)    <= sub_wire92(14);
	sub_wire1(36, 15)    <= sub_wire92(15);
	sub_wire1(36, 16)    <= sub_wire92(16);
	sub_wire1(36, 17)    <= sub_wire92(17);
	sub_wire1(36, 18)    <= sub_wire92(18);
	sub_wire1(36, 19)    <= sub_wire92(19);
	sub_wire1(36, 20)    <= sub_wire92(20);
	sub_wire1(36, 21)    <= sub_wire92(21);
	sub_wire1(36, 22)    <= sub_wire92(22);
	sub_wire1(36, 23)    <= sub_wire92(23);
	sub_wire1(36, 24)    <= sub_wire92(24);
	sub_wire1(36, 25)    <= sub_wire92(25);
	sub_wire1(36, 26)    <= sub_wire92(26);
	sub_wire1(36, 27)    <= sub_wire92(27);
	sub_wire1(36, 28)    <= sub_wire92(28);
	sub_wire1(36, 29)    <= sub_wire92(29);
	sub_wire1(36, 30)    <= sub_wire92(30);
	sub_wire1(36, 31)    <= sub_wire92(31);
	sub_wire1(35, 0)    <= sub_wire93(0);
	sub_wire1(35, 1)    <= sub_wire93(1);
	sub_wire1(35, 2)    <= sub_wire93(2);
	sub_wire1(35, 3)    <= sub_wire93(3);
	sub_wire1(35, 4)    <= sub_wire93(4);
	sub_wire1(35, 5)    <= sub_wire93(5);
	sub_wire1(35, 6)    <= sub_wire93(6);
	sub_wire1(35, 7)    <= sub_wire93(7);
	sub_wire1(35, 8)    <= sub_wire93(8);
	sub_wire1(35, 9)    <= sub_wire93(9);
	sub_wire1(35, 10)    <= sub_wire93(10);
	sub_wire1(35, 11)    <= sub_wire93(11);
	sub_wire1(35, 12)    <= sub_wire93(12);
	sub_wire1(35, 13)    <= sub_wire93(13);
	sub_wire1(35, 14)    <= sub_wire93(14);
	sub_wire1(35, 15)    <= sub_wire93(15);
	sub_wire1(35, 16)    <= sub_wire93(16);
	sub_wire1(35, 17)    <= sub_wire93(17);
	sub_wire1(35, 18)    <= sub_wire93(18);
	sub_wire1(35, 19)    <= sub_wire93(19);
	sub_wire1(35, 20)    <= sub_wire93(20);
	sub_wire1(35, 21)    <= sub_wire93(21);
	sub_wire1(35, 22)    <= sub_wire93(22);
	sub_wire1(35, 23)    <= sub_wire93(23);
	sub_wire1(35, 24)    <= sub_wire93(24);
	sub_wire1(35, 25)    <= sub_wire93(25);
	sub_wire1(35, 26)    <= sub_wire93(26);
	sub_wire1(35, 27)    <= sub_wire93(27);
	sub_wire1(35, 28)    <= sub_wire93(28);
	sub_wire1(35, 29)    <= sub_wire93(29);
	sub_wire1(35, 30)    <= sub_wire93(30);
	sub_wire1(35, 31)    <= sub_wire93(31);
	sub_wire1(34, 0)    <= sub_wire94(0);
	sub_wire1(34, 1)    <= sub_wire94(1);
	sub_wire1(34, 2)    <= sub_wire94(2);
	sub_wire1(34, 3)    <= sub_wire94(3);
	sub_wire1(34, 4)    <= sub_wire94(4);
	sub_wire1(34, 5)    <= sub_wire94(5);
	sub_wire1(34, 6)    <= sub_wire94(6);
	sub_wire1(34, 7)    <= sub_wire94(7);
	sub_wire1(34, 8)    <= sub_wire94(8);
	sub_wire1(34, 9)    <= sub_wire94(9);
	sub_wire1(34, 10)    <= sub_wire94(10);
	sub_wire1(34, 11)    <= sub_wire94(11);
	sub_wire1(34, 12)    <= sub_wire94(12);
	sub_wire1(34, 13)    <= sub_wire94(13);
	sub_wire1(34, 14)    <= sub_wire94(14);
	sub_wire1(34, 15)    <= sub_wire94(15);
	sub_wire1(34, 16)    <= sub_wire94(16);
	sub_wire1(34, 17)    <= sub_wire94(17);
	sub_wire1(34, 18)    <= sub_wire94(18);
	sub_wire1(34, 19)    <= sub_wire94(19);
	sub_wire1(34, 20)    <= sub_wire94(20);
	sub_wire1(34, 21)    <= sub_wire94(21);
	sub_wire1(34, 22)    <= sub_wire94(22);
	sub_wire1(34, 23)    <= sub_wire94(23);
	sub_wire1(34, 24)    <= sub_wire94(24);
	sub_wire1(34, 25)    <= sub_wire94(25);
	sub_wire1(34, 26)    <= sub_wire94(26);
	sub_wire1(34, 27)    <= sub_wire94(27);
	sub_wire1(34, 28)    <= sub_wire94(28);
	sub_wire1(34, 29)    <= sub_wire94(29);
	sub_wire1(34, 30)    <= sub_wire94(30);
	sub_wire1(34, 31)    <= sub_wire94(31);
	sub_wire1(33, 0)    <= sub_wire95(0);
	sub_wire1(33, 1)    <= sub_wire95(1);
	sub_wire1(33, 2)    <= sub_wire95(2);
	sub_wire1(33, 3)    <= sub_wire95(3);
	sub_wire1(33, 4)    <= sub_wire95(4);
	sub_wire1(33, 5)    <= sub_wire95(5);
	sub_wire1(33, 6)    <= sub_wire95(6);
	sub_wire1(33, 7)    <= sub_wire95(7);
	sub_wire1(33, 8)    <= sub_wire95(8);
	sub_wire1(33, 9)    <= sub_wire95(9);
	sub_wire1(33, 10)    <= sub_wire95(10);
	sub_wire1(33, 11)    <= sub_wire95(11);
	sub_wire1(33, 12)    <= sub_wire95(12);
	sub_wire1(33, 13)    <= sub_wire95(13);
	sub_wire1(33, 14)    <= sub_wire95(14);
	sub_wire1(33, 15)    <= sub_wire95(15);
	sub_wire1(33, 16)    <= sub_wire95(16);
	sub_wire1(33, 17)    <= sub_wire95(17);
	sub_wire1(33, 18)    <= sub_wire95(18);
	sub_wire1(33, 19)    <= sub_wire95(19);
	sub_wire1(33, 20)    <= sub_wire95(20);
	sub_wire1(33, 21)    <= sub_wire95(21);
	sub_wire1(33, 22)    <= sub_wire95(22);
	sub_wire1(33, 23)    <= sub_wire95(23);
	sub_wire1(33, 24)    <= sub_wire95(24);
	sub_wire1(33, 25)    <= sub_wire95(25);
	sub_wire1(33, 26)    <= sub_wire95(26);
	sub_wire1(33, 27)    <= sub_wire95(27);
	sub_wire1(33, 28)    <= sub_wire95(28);
	sub_wire1(33, 29)    <= sub_wire95(29);
	sub_wire1(33, 30)    <= sub_wire95(30);
	sub_wire1(33, 31)    <= sub_wire95(31);
	sub_wire1(32, 0)    <= sub_wire96(0);
	sub_wire1(32, 1)    <= sub_wire96(1);
	sub_wire1(32, 2)    <= sub_wire96(2);
	sub_wire1(32, 3)    <= sub_wire96(3);
	sub_wire1(32, 4)    <= sub_wire96(4);
	sub_wire1(32, 5)    <= sub_wire96(5);
	sub_wire1(32, 6)    <= sub_wire96(6);
	sub_wire1(32, 7)    <= sub_wire96(7);
	sub_wire1(32, 8)    <= sub_wire96(8);
	sub_wire1(32, 9)    <= sub_wire96(9);
	sub_wire1(32, 10)    <= sub_wire96(10);
	sub_wire1(32, 11)    <= sub_wire96(11);
	sub_wire1(32, 12)    <= sub_wire96(12);
	sub_wire1(32, 13)    <= sub_wire96(13);
	sub_wire1(32, 14)    <= sub_wire96(14);
	sub_wire1(32, 15)    <= sub_wire96(15);
	sub_wire1(32, 16)    <= sub_wire96(16);
	sub_wire1(32, 17)    <= sub_wire96(17);
	sub_wire1(32, 18)    <= sub_wire96(18);
	sub_wire1(32, 19)    <= sub_wire96(19);
	sub_wire1(32, 20)    <= sub_wire96(20);
	sub_wire1(32, 21)    <= sub_wire96(21);
	sub_wire1(32, 22)    <= sub_wire96(22);
	sub_wire1(32, 23)    <= sub_wire96(23);
	sub_wire1(32, 24)    <= sub_wire96(24);
	sub_wire1(32, 25)    <= sub_wire96(25);
	sub_wire1(32, 26)    <= sub_wire96(26);
	sub_wire1(32, 27)    <= sub_wire96(27);
	sub_wire1(32, 28)    <= sub_wire96(28);
	sub_wire1(32, 29)    <= sub_wire96(29);
	sub_wire1(32, 30)    <= sub_wire96(30);
	sub_wire1(32, 31)    <= sub_wire96(31);
	sub_wire1(31, 0)    <= sub_wire97(0);
	sub_wire1(31, 1)    <= sub_wire97(1);
	sub_wire1(31, 2)    <= sub_wire97(2);
	sub_wire1(31, 3)    <= sub_wire97(3);
	sub_wire1(31, 4)    <= sub_wire97(4);
	sub_wire1(31, 5)    <= sub_wire97(5);
	sub_wire1(31, 6)    <= sub_wire97(6);
	sub_wire1(31, 7)    <= sub_wire97(7);
	sub_wire1(31, 8)    <= sub_wire97(8);
	sub_wire1(31, 9)    <= sub_wire97(9);
	sub_wire1(31, 10)    <= sub_wire97(10);
	sub_wire1(31, 11)    <= sub_wire97(11);
	sub_wire1(31, 12)    <= sub_wire97(12);
	sub_wire1(31, 13)    <= sub_wire97(13);
	sub_wire1(31, 14)    <= sub_wire97(14);
	sub_wire1(31, 15)    <= sub_wire97(15);
	sub_wire1(31, 16)    <= sub_wire97(16);
	sub_wire1(31, 17)    <= sub_wire97(17);
	sub_wire1(31, 18)    <= sub_wire97(18);
	sub_wire1(31, 19)    <= sub_wire97(19);
	sub_wire1(31, 20)    <= sub_wire97(20);
	sub_wire1(31, 21)    <= sub_wire97(21);
	sub_wire1(31, 22)    <= sub_wire97(22);
	sub_wire1(31, 23)    <= sub_wire97(23);
	sub_wire1(31, 24)    <= sub_wire97(24);
	sub_wire1(31, 25)    <= sub_wire97(25);
	sub_wire1(31, 26)    <= sub_wire97(26);
	sub_wire1(31, 27)    <= sub_wire97(27);
	sub_wire1(31, 28)    <= sub_wire97(28);
	sub_wire1(31, 29)    <= sub_wire97(29);
	sub_wire1(31, 30)    <= sub_wire97(30);
	sub_wire1(31, 31)    <= sub_wire97(31);
	sub_wire1(30, 0)    <= sub_wire98(0);
	sub_wire1(30, 1)    <= sub_wire98(1);
	sub_wire1(30, 2)    <= sub_wire98(2);
	sub_wire1(30, 3)    <= sub_wire98(3);
	sub_wire1(30, 4)    <= sub_wire98(4);
	sub_wire1(30, 5)    <= sub_wire98(5);
	sub_wire1(30, 6)    <= sub_wire98(6);
	sub_wire1(30, 7)    <= sub_wire98(7);
	sub_wire1(30, 8)    <= sub_wire98(8);
	sub_wire1(30, 9)    <= sub_wire98(9);
	sub_wire1(30, 10)    <= sub_wire98(10);
	sub_wire1(30, 11)    <= sub_wire98(11);
	sub_wire1(30, 12)    <= sub_wire98(12);
	sub_wire1(30, 13)    <= sub_wire98(13);
	sub_wire1(30, 14)    <= sub_wire98(14);
	sub_wire1(30, 15)    <= sub_wire98(15);
	sub_wire1(30, 16)    <= sub_wire98(16);
	sub_wire1(30, 17)    <= sub_wire98(17);
	sub_wire1(30, 18)    <= sub_wire98(18);
	sub_wire1(30, 19)    <= sub_wire98(19);
	sub_wire1(30, 20)    <= sub_wire98(20);
	sub_wire1(30, 21)    <= sub_wire98(21);
	sub_wire1(30, 22)    <= sub_wire98(22);
	sub_wire1(30, 23)    <= sub_wire98(23);
	sub_wire1(30, 24)    <= sub_wire98(24);
	sub_wire1(30, 25)    <= sub_wire98(25);
	sub_wire1(30, 26)    <= sub_wire98(26);
	sub_wire1(30, 27)    <= sub_wire98(27);
	sub_wire1(30, 28)    <= sub_wire98(28);
	sub_wire1(30, 29)    <= sub_wire98(29);
	sub_wire1(30, 30)    <= sub_wire98(30);
	sub_wire1(30, 31)    <= sub_wire98(31);
	sub_wire1(29, 0)    <= sub_wire99(0);
	sub_wire1(29, 1)    <= sub_wire99(1);
	sub_wire1(29, 2)    <= sub_wire99(2);
	sub_wire1(29, 3)    <= sub_wire99(3);
	sub_wire1(29, 4)    <= sub_wire99(4);
	sub_wire1(29, 5)    <= sub_wire99(5);
	sub_wire1(29, 6)    <= sub_wire99(6);
	sub_wire1(29, 7)    <= sub_wire99(7);
	sub_wire1(29, 8)    <= sub_wire99(8);
	sub_wire1(29, 9)    <= sub_wire99(9);
	sub_wire1(29, 10)    <= sub_wire99(10);
	sub_wire1(29, 11)    <= sub_wire99(11);
	sub_wire1(29, 12)    <= sub_wire99(12);
	sub_wire1(29, 13)    <= sub_wire99(13);
	sub_wire1(29, 14)    <= sub_wire99(14);
	sub_wire1(29, 15)    <= sub_wire99(15);
	sub_wire1(29, 16)    <= sub_wire99(16);
	sub_wire1(29, 17)    <= sub_wire99(17);
	sub_wire1(29, 18)    <= sub_wire99(18);
	sub_wire1(29, 19)    <= sub_wire99(19);
	sub_wire1(29, 20)    <= sub_wire99(20);
	sub_wire1(29, 21)    <= sub_wire99(21);
	sub_wire1(29, 22)    <= sub_wire99(22);
	sub_wire1(29, 23)    <= sub_wire99(23);
	sub_wire1(29, 24)    <= sub_wire99(24);
	sub_wire1(29, 25)    <= sub_wire99(25);
	sub_wire1(29, 26)    <= sub_wire99(26);
	sub_wire1(29, 27)    <= sub_wire99(27);
	sub_wire1(29, 28)    <= sub_wire99(28);
	sub_wire1(29, 29)    <= sub_wire99(29);
	sub_wire1(29, 30)    <= sub_wire99(30);
	sub_wire1(29, 31)    <= sub_wire99(31);
	sub_wire1(28, 0)    <= sub_wire100(0);
	sub_wire1(28, 1)    <= sub_wire100(1);
	sub_wire1(28, 2)    <= sub_wire100(2);
	sub_wire1(28, 3)    <= sub_wire100(3);
	sub_wire1(28, 4)    <= sub_wire100(4);
	sub_wire1(28, 5)    <= sub_wire100(5);
	sub_wire1(28, 6)    <= sub_wire100(6);
	sub_wire1(28, 7)    <= sub_wire100(7);
	sub_wire1(28, 8)    <= sub_wire100(8);
	sub_wire1(28, 9)    <= sub_wire100(9);
	sub_wire1(28, 10)    <= sub_wire100(10);
	sub_wire1(28, 11)    <= sub_wire100(11);
	sub_wire1(28, 12)    <= sub_wire100(12);
	sub_wire1(28, 13)    <= sub_wire100(13);
	sub_wire1(28, 14)    <= sub_wire100(14);
	sub_wire1(28, 15)    <= sub_wire100(15);
	sub_wire1(28, 16)    <= sub_wire100(16);
	sub_wire1(28, 17)    <= sub_wire100(17);
	sub_wire1(28, 18)    <= sub_wire100(18);
	sub_wire1(28, 19)    <= sub_wire100(19);
	sub_wire1(28, 20)    <= sub_wire100(20);
	sub_wire1(28, 21)    <= sub_wire100(21);
	sub_wire1(28, 22)    <= sub_wire100(22);
	sub_wire1(28, 23)    <= sub_wire100(23);
	sub_wire1(28, 24)    <= sub_wire100(24);
	sub_wire1(28, 25)    <= sub_wire100(25);
	sub_wire1(28, 26)    <= sub_wire100(26);
	sub_wire1(28, 27)    <= sub_wire100(27);
	sub_wire1(28, 28)    <= sub_wire100(28);
	sub_wire1(28, 29)    <= sub_wire100(29);
	sub_wire1(28, 30)    <= sub_wire100(30);
	sub_wire1(28, 31)    <= sub_wire100(31);
	sub_wire1(27, 0)    <= sub_wire101(0);
	sub_wire1(27, 1)    <= sub_wire101(1);
	sub_wire1(27, 2)    <= sub_wire101(2);
	sub_wire1(27, 3)    <= sub_wire101(3);
	sub_wire1(27, 4)    <= sub_wire101(4);
	sub_wire1(27, 5)    <= sub_wire101(5);
	sub_wire1(27, 6)    <= sub_wire101(6);
	sub_wire1(27, 7)    <= sub_wire101(7);
	sub_wire1(27, 8)    <= sub_wire101(8);
	sub_wire1(27, 9)    <= sub_wire101(9);
	sub_wire1(27, 10)    <= sub_wire101(10);
	sub_wire1(27, 11)    <= sub_wire101(11);
	sub_wire1(27, 12)    <= sub_wire101(12);
	sub_wire1(27, 13)    <= sub_wire101(13);
	sub_wire1(27, 14)    <= sub_wire101(14);
	sub_wire1(27, 15)    <= sub_wire101(15);
	sub_wire1(27, 16)    <= sub_wire101(16);
	sub_wire1(27, 17)    <= sub_wire101(17);
	sub_wire1(27, 18)    <= sub_wire101(18);
	sub_wire1(27, 19)    <= sub_wire101(19);
	sub_wire1(27, 20)    <= sub_wire101(20);
	sub_wire1(27, 21)    <= sub_wire101(21);
	sub_wire1(27, 22)    <= sub_wire101(22);
	sub_wire1(27, 23)    <= sub_wire101(23);
	sub_wire1(27, 24)    <= sub_wire101(24);
	sub_wire1(27, 25)    <= sub_wire101(25);
	sub_wire1(27, 26)    <= sub_wire101(26);
	sub_wire1(27, 27)    <= sub_wire101(27);
	sub_wire1(27, 28)    <= sub_wire101(28);
	sub_wire1(27, 29)    <= sub_wire101(29);
	sub_wire1(27, 30)    <= sub_wire101(30);
	sub_wire1(27, 31)    <= sub_wire101(31);
	sub_wire1(26, 0)    <= sub_wire102(0);
	sub_wire1(26, 1)    <= sub_wire102(1);
	sub_wire1(26, 2)    <= sub_wire102(2);
	sub_wire1(26, 3)    <= sub_wire102(3);
	sub_wire1(26, 4)    <= sub_wire102(4);
	sub_wire1(26, 5)    <= sub_wire102(5);
	sub_wire1(26, 6)    <= sub_wire102(6);
	sub_wire1(26, 7)    <= sub_wire102(7);
	sub_wire1(26, 8)    <= sub_wire102(8);
	sub_wire1(26, 9)    <= sub_wire102(9);
	sub_wire1(26, 10)    <= sub_wire102(10);
	sub_wire1(26, 11)    <= sub_wire102(11);
	sub_wire1(26, 12)    <= sub_wire102(12);
	sub_wire1(26, 13)    <= sub_wire102(13);
	sub_wire1(26, 14)    <= sub_wire102(14);
	sub_wire1(26, 15)    <= sub_wire102(15);
	sub_wire1(26, 16)    <= sub_wire102(16);
	sub_wire1(26, 17)    <= sub_wire102(17);
	sub_wire1(26, 18)    <= sub_wire102(18);
	sub_wire1(26, 19)    <= sub_wire102(19);
	sub_wire1(26, 20)    <= sub_wire102(20);
	sub_wire1(26, 21)    <= sub_wire102(21);
	sub_wire1(26, 22)    <= sub_wire102(22);
	sub_wire1(26, 23)    <= sub_wire102(23);
	sub_wire1(26, 24)    <= sub_wire102(24);
	sub_wire1(26, 25)    <= sub_wire102(25);
	sub_wire1(26, 26)    <= sub_wire102(26);
	sub_wire1(26, 27)    <= sub_wire102(27);
	sub_wire1(26, 28)    <= sub_wire102(28);
	sub_wire1(26, 29)    <= sub_wire102(29);
	sub_wire1(26, 30)    <= sub_wire102(30);
	sub_wire1(26, 31)    <= sub_wire102(31);
	sub_wire1(25, 0)    <= sub_wire103(0);
	sub_wire1(25, 1)    <= sub_wire103(1);
	sub_wire1(25, 2)    <= sub_wire103(2);
	sub_wire1(25, 3)    <= sub_wire103(3);
	sub_wire1(25, 4)    <= sub_wire103(4);
	sub_wire1(25, 5)    <= sub_wire103(5);
	sub_wire1(25, 6)    <= sub_wire103(6);
	sub_wire1(25, 7)    <= sub_wire103(7);
	sub_wire1(25, 8)    <= sub_wire103(8);
	sub_wire1(25, 9)    <= sub_wire103(9);
	sub_wire1(25, 10)    <= sub_wire103(10);
	sub_wire1(25, 11)    <= sub_wire103(11);
	sub_wire1(25, 12)    <= sub_wire103(12);
	sub_wire1(25, 13)    <= sub_wire103(13);
	sub_wire1(25, 14)    <= sub_wire103(14);
	sub_wire1(25, 15)    <= sub_wire103(15);
	sub_wire1(25, 16)    <= sub_wire103(16);
	sub_wire1(25, 17)    <= sub_wire103(17);
	sub_wire1(25, 18)    <= sub_wire103(18);
	sub_wire1(25, 19)    <= sub_wire103(19);
	sub_wire1(25, 20)    <= sub_wire103(20);
	sub_wire1(25, 21)    <= sub_wire103(21);
	sub_wire1(25, 22)    <= sub_wire103(22);
	sub_wire1(25, 23)    <= sub_wire103(23);
	sub_wire1(25, 24)    <= sub_wire103(24);
	sub_wire1(25, 25)    <= sub_wire103(25);
	sub_wire1(25, 26)    <= sub_wire103(26);
	sub_wire1(25, 27)    <= sub_wire103(27);
	sub_wire1(25, 28)    <= sub_wire103(28);
	sub_wire1(25, 29)    <= sub_wire103(29);
	sub_wire1(25, 30)    <= sub_wire103(30);
	sub_wire1(25, 31)    <= sub_wire103(31);
	sub_wire1(24, 0)    <= sub_wire104(0);
	sub_wire1(24, 1)    <= sub_wire104(1);
	sub_wire1(24, 2)    <= sub_wire104(2);
	sub_wire1(24, 3)    <= sub_wire104(3);
	sub_wire1(24, 4)    <= sub_wire104(4);
	sub_wire1(24, 5)    <= sub_wire104(5);
	sub_wire1(24, 6)    <= sub_wire104(6);
	sub_wire1(24, 7)    <= sub_wire104(7);
	sub_wire1(24, 8)    <= sub_wire104(8);
	sub_wire1(24, 9)    <= sub_wire104(9);
	sub_wire1(24, 10)    <= sub_wire104(10);
	sub_wire1(24, 11)    <= sub_wire104(11);
	sub_wire1(24, 12)    <= sub_wire104(12);
	sub_wire1(24, 13)    <= sub_wire104(13);
	sub_wire1(24, 14)    <= sub_wire104(14);
	sub_wire1(24, 15)    <= sub_wire104(15);
	sub_wire1(24, 16)    <= sub_wire104(16);
	sub_wire1(24, 17)    <= sub_wire104(17);
	sub_wire1(24, 18)    <= sub_wire104(18);
	sub_wire1(24, 19)    <= sub_wire104(19);
	sub_wire1(24, 20)    <= sub_wire104(20);
	sub_wire1(24, 21)    <= sub_wire104(21);
	sub_wire1(24, 22)    <= sub_wire104(22);
	sub_wire1(24, 23)    <= sub_wire104(23);
	sub_wire1(24, 24)    <= sub_wire104(24);
	sub_wire1(24, 25)    <= sub_wire104(25);
	sub_wire1(24, 26)    <= sub_wire104(26);
	sub_wire1(24, 27)    <= sub_wire104(27);
	sub_wire1(24, 28)    <= sub_wire104(28);
	sub_wire1(24, 29)    <= sub_wire104(29);
	sub_wire1(24, 30)    <= sub_wire104(30);
	sub_wire1(24, 31)    <= sub_wire104(31);
	sub_wire1(23, 0)    <= sub_wire105(0);
	sub_wire1(23, 1)    <= sub_wire105(1);
	sub_wire1(23, 2)    <= sub_wire105(2);
	sub_wire1(23, 3)    <= sub_wire105(3);
	sub_wire1(23, 4)    <= sub_wire105(4);
	sub_wire1(23, 5)    <= sub_wire105(5);
	sub_wire1(23, 6)    <= sub_wire105(6);
	sub_wire1(23, 7)    <= sub_wire105(7);
	sub_wire1(23, 8)    <= sub_wire105(8);
	sub_wire1(23, 9)    <= sub_wire105(9);
	sub_wire1(23, 10)    <= sub_wire105(10);
	sub_wire1(23, 11)    <= sub_wire105(11);
	sub_wire1(23, 12)    <= sub_wire105(12);
	sub_wire1(23, 13)    <= sub_wire105(13);
	sub_wire1(23, 14)    <= sub_wire105(14);
	sub_wire1(23, 15)    <= sub_wire105(15);
	sub_wire1(23, 16)    <= sub_wire105(16);
	sub_wire1(23, 17)    <= sub_wire105(17);
	sub_wire1(23, 18)    <= sub_wire105(18);
	sub_wire1(23, 19)    <= sub_wire105(19);
	sub_wire1(23, 20)    <= sub_wire105(20);
	sub_wire1(23, 21)    <= sub_wire105(21);
	sub_wire1(23, 22)    <= sub_wire105(22);
	sub_wire1(23, 23)    <= sub_wire105(23);
	sub_wire1(23, 24)    <= sub_wire105(24);
	sub_wire1(23, 25)    <= sub_wire105(25);
	sub_wire1(23, 26)    <= sub_wire105(26);
	sub_wire1(23, 27)    <= sub_wire105(27);
	sub_wire1(23, 28)    <= sub_wire105(28);
	sub_wire1(23, 29)    <= sub_wire105(29);
	sub_wire1(23, 30)    <= sub_wire105(30);
	sub_wire1(23, 31)    <= sub_wire105(31);
	sub_wire1(22, 0)    <= sub_wire106(0);
	sub_wire1(22, 1)    <= sub_wire106(1);
	sub_wire1(22, 2)    <= sub_wire106(2);
	sub_wire1(22, 3)    <= sub_wire106(3);
	sub_wire1(22, 4)    <= sub_wire106(4);
	sub_wire1(22, 5)    <= sub_wire106(5);
	sub_wire1(22, 6)    <= sub_wire106(6);
	sub_wire1(22, 7)    <= sub_wire106(7);
	sub_wire1(22, 8)    <= sub_wire106(8);
	sub_wire1(22, 9)    <= sub_wire106(9);
	sub_wire1(22, 10)    <= sub_wire106(10);
	sub_wire1(22, 11)    <= sub_wire106(11);
	sub_wire1(22, 12)    <= sub_wire106(12);
	sub_wire1(22, 13)    <= sub_wire106(13);
	sub_wire1(22, 14)    <= sub_wire106(14);
	sub_wire1(22, 15)    <= sub_wire106(15);
	sub_wire1(22, 16)    <= sub_wire106(16);
	sub_wire1(22, 17)    <= sub_wire106(17);
	sub_wire1(22, 18)    <= sub_wire106(18);
	sub_wire1(22, 19)    <= sub_wire106(19);
	sub_wire1(22, 20)    <= sub_wire106(20);
	sub_wire1(22, 21)    <= sub_wire106(21);
	sub_wire1(22, 22)    <= sub_wire106(22);
	sub_wire1(22, 23)    <= sub_wire106(23);
	sub_wire1(22, 24)    <= sub_wire106(24);
	sub_wire1(22, 25)    <= sub_wire106(25);
	sub_wire1(22, 26)    <= sub_wire106(26);
	sub_wire1(22, 27)    <= sub_wire106(27);
	sub_wire1(22, 28)    <= sub_wire106(28);
	sub_wire1(22, 29)    <= sub_wire106(29);
	sub_wire1(22, 30)    <= sub_wire106(30);
	sub_wire1(22, 31)    <= sub_wire106(31);
	sub_wire1(21, 0)    <= sub_wire107(0);
	sub_wire1(21, 1)    <= sub_wire107(1);
	sub_wire1(21, 2)    <= sub_wire107(2);
	sub_wire1(21, 3)    <= sub_wire107(3);
	sub_wire1(21, 4)    <= sub_wire107(4);
	sub_wire1(21, 5)    <= sub_wire107(5);
	sub_wire1(21, 6)    <= sub_wire107(6);
	sub_wire1(21, 7)    <= sub_wire107(7);
	sub_wire1(21, 8)    <= sub_wire107(8);
	sub_wire1(21, 9)    <= sub_wire107(9);
	sub_wire1(21, 10)    <= sub_wire107(10);
	sub_wire1(21, 11)    <= sub_wire107(11);
	sub_wire1(21, 12)    <= sub_wire107(12);
	sub_wire1(21, 13)    <= sub_wire107(13);
	sub_wire1(21, 14)    <= sub_wire107(14);
	sub_wire1(21, 15)    <= sub_wire107(15);
	sub_wire1(21, 16)    <= sub_wire107(16);
	sub_wire1(21, 17)    <= sub_wire107(17);
	sub_wire1(21, 18)    <= sub_wire107(18);
	sub_wire1(21, 19)    <= sub_wire107(19);
	sub_wire1(21, 20)    <= sub_wire107(20);
	sub_wire1(21, 21)    <= sub_wire107(21);
	sub_wire1(21, 22)    <= sub_wire107(22);
	sub_wire1(21, 23)    <= sub_wire107(23);
	sub_wire1(21, 24)    <= sub_wire107(24);
	sub_wire1(21, 25)    <= sub_wire107(25);
	sub_wire1(21, 26)    <= sub_wire107(26);
	sub_wire1(21, 27)    <= sub_wire107(27);
	sub_wire1(21, 28)    <= sub_wire107(28);
	sub_wire1(21, 29)    <= sub_wire107(29);
	sub_wire1(21, 30)    <= sub_wire107(30);
	sub_wire1(21, 31)    <= sub_wire107(31);
	sub_wire1(20, 0)    <= sub_wire108(0);
	sub_wire1(20, 1)    <= sub_wire108(1);
	sub_wire1(20, 2)    <= sub_wire108(2);
	sub_wire1(20, 3)    <= sub_wire108(3);
	sub_wire1(20, 4)    <= sub_wire108(4);
	sub_wire1(20, 5)    <= sub_wire108(5);
	sub_wire1(20, 6)    <= sub_wire108(6);
	sub_wire1(20, 7)    <= sub_wire108(7);
	sub_wire1(20, 8)    <= sub_wire108(8);
	sub_wire1(20, 9)    <= sub_wire108(9);
	sub_wire1(20, 10)    <= sub_wire108(10);
	sub_wire1(20, 11)    <= sub_wire108(11);
	sub_wire1(20, 12)    <= sub_wire108(12);
	sub_wire1(20, 13)    <= sub_wire108(13);
	sub_wire1(20, 14)    <= sub_wire108(14);
	sub_wire1(20, 15)    <= sub_wire108(15);
	sub_wire1(20, 16)    <= sub_wire108(16);
	sub_wire1(20, 17)    <= sub_wire108(17);
	sub_wire1(20, 18)    <= sub_wire108(18);
	sub_wire1(20, 19)    <= sub_wire108(19);
	sub_wire1(20, 20)    <= sub_wire108(20);
	sub_wire1(20, 21)    <= sub_wire108(21);
	sub_wire1(20, 22)    <= sub_wire108(22);
	sub_wire1(20, 23)    <= sub_wire108(23);
	sub_wire1(20, 24)    <= sub_wire108(24);
	sub_wire1(20, 25)    <= sub_wire108(25);
	sub_wire1(20, 26)    <= sub_wire108(26);
	sub_wire1(20, 27)    <= sub_wire108(27);
	sub_wire1(20, 28)    <= sub_wire108(28);
	sub_wire1(20, 29)    <= sub_wire108(29);
	sub_wire1(20, 30)    <= sub_wire108(30);
	sub_wire1(20, 31)    <= sub_wire108(31);
	sub_wire1(19, 0)    <= sub_wire109(0);
	sub_wire1(19, 1)    <= sub_wire109(1);
	sub_wire1(19, 2)    <= sub_wire109(2);
	sub_wire1(19, 3)    <= sub_wire109(3);
	sub_wire1(19, 4)    <= sub_wire109(4);
	sub_wire1(19, 5)    <= sub_wire109(5);
	sub_wire1(19, 6)    <= sub_wire109(6);
	sub_wire1(19, 7)    <= sub_wire109(7);
	sub_wire1(19, 8)    <= sub_wire109(8);
	sub_wire1(19, 9)    <= sub_wire109(9);
	sub_wire1(19, 10)    <= sub_wire109(10);
	sub_wire1(19, 11)    <= sub_wire109(11);
	sub_wire1(19, 12)    <= sub_wire109(12);
	sub_wire1(19, 13)    <= sub_wire109(13);
	sub_wire1(19, 14)    <= sub_wire109(14);
	sub_wire1(19, 15)    <= sub_wire109(15);
	sub_wire1(19, 16)    <= sub_wire109(16);
	sub_wire1(19, 17)    <= sub_wire109(17);
	sub_wire1(19, 18)    <= sub_wire109(18);
	sub_wire1(19, 19)    <= sub_wire109(19);
	sub_wire1(19, 20)    <= sub_wire109(20);
	sub_wire1(19, 21)    <= sub_wire109(21);
	sub_wire1(19, 22)    <= sub_wire109(22);
	sub_wire1(19, 23)    <= sub_wire109(23);
	sub_wire1(19, 24)    <= sub_wire109(24);
	sub_wire1(19, 25)    <= sub_wire109(25);
	sub_wire1(19, 26)    <= sub_wire109(26);
	sub_wire1(19, 27)    <= sub_wire109(27);
	sub_wire1(19, 28)    <= sub_wire109(28);
	sub_wire1(19, 29)    <= sub_wire109(29);
	sub_wire1(19, 30)    <= sub_wire109(30);
	sub_wire1(19, 31)    <= sub_wire109(31);
	sub_wire1(18, 0)    <= sub_wire110(0);
	sub_wire1(18, 1)    <= sub_wire110(1);
	sub_wire1(18, 2)    <= sub_wire110(2);
	sub_wire1(18, 3)    <= sub_wire110(3);
	sub_wire1(18, 4)    <= sub_wire110(4);
	sub_wire1(18, 5)    <= sub_wire110(5);
	sub_wire1(18, 6)    <= sub_wire110(6);
	sub_wire1(18, 7)    <= sub_wire110(7);
	sub_wire1(18, 8)    <= sub_wire110(8);
	sub_wire1(18, 9)    <= sub_wire110(9);
	sub_wire1(18, 10)    <= sub_wire110(10);
	sub_wire1(18, 11)    <= sub_wire110(11);
	sub_wire1(18, 12)    <= sub_wire110(12);
	sub_wire1(18, 13)    <= sub_wire110(13);
	sub_wire1(18, 14)    <= sub_wire110(14);
	sub_wire1(18, 15)    <= sub_wire110(15);
	sub_wire1(18, 16)    <= sub_wire110(16);
	sub_wire1(18, 17)    <= sub_wire110(17);
	sub_wire1(18, 18)    <= sub_wire110(18);
	sub_wire1(18, 19)    <= sub_wire110(19);
	sub_wire1(18, 20)    <= sub_wire110(20);
	sub_wire1(18, 21)    <= sub_wire110(21);
	sub_wire1(18, 22)    <= sub_wire110(22);
	sub_wire1(18, 23)    <= sub_wire110(23);
	sub_wire1(18, 24)    <= sub_wire110(24);
	sub_wire1(18, 25)    <= sub_wire110(25);
	sub_wire1(18, 26)    <= sub_wire110(26);
	sub_wire1(18, 27)    <= sub_wire110(27);
	sub_wire1(18, 28)    <= sub_wire110(28);
	sub_wire1(18, 29)    <= sub_wire110(29);
	sub_wire1(18, 30)    <= sub_wire110(30);
	sub_wire1(18, 31)    <= sub_wire110(31);
	sub_wire1(17, 0)    <= sub_wire111(0);
	sub_wire1(17, 1)    <= sub_wire111(1);
	sub_wire1(17, 2)    <= sub_wire111(2);
	sub_wire1(17, 3)    <= sub_wire111(3);
	sub_wire1(17, 4)    <= sub_wire111(4);
	sub_wire1(17, 5)    <= sub_wire111(5);
	sub_wire1(17, 6)    <= sub_wire111(6);
	sub_wire1(17, 7)    <= sub_wire111(7);
	sub_wire1(17, 8)    <= sub_wire111(8);
	sub_wire1(17, 9)    <= sub_wire111(9);
	sub_wire1(17, 10)    <= sub_wire111(10);
	sub_wire1(17, 11)    <= sub_wire111(11);
	sub_wire1(17, 12)    <= sub_wire111(12);
	sub_wire1(17, 13)    <= sub_wire111(13);
	sub_wire1(17, 14)    <= sub_wire111(14);
	sub_wire1(17, 15)    <= sub_wire111(15);
	sub_wire1(17, 16)    <= sub_wire111(16);
	sub_wire1(17, 17)    <= sub_wire111(17);
	sub_wire1(17, 18)    <= sub_wire111(18);
	sub_wire1(17, 19)    <= sub_wire111(19);
	sub_wire1(17, 20)    <= sub_wire111(20);
	sub_wire1(17, 21)    <= sub_wire111(21);
	sub_wire1(17, 22)    <= sub_wire111(22);
	sub_wire1(17, 23)    <= sub_wire111(23);
	sub_wire1(17, 24)    <= sub_wire111(24);
	sub_wire1(17, 25)    <= sub_wire111(25);
	sub_wire1(17, 26)    <= sub_wire111(26);
	sub_wire1(17, 27)    <= sub_wire111(27);
	sub_wire1(17, 28)    <= sub_wire111(28);
	sub_wire1(17, 29)    <= sub_wire111(29);
	sub_wire1(17, 30)    <= sub_wire111(30);
	sub_wire1(17, 31)    <= sub_wire111(31);
	sub_wire1(16, 0)    <= sub_wire112(0);
	sub_wire1(16, 1)    <= sub_wire112(1);
	sub_wire1(16, 2)    <= sub_wire112(2);
	sub_wire1(16, 3)    <= sub_wire112(3);
	sub_wire1(16, 4)    <= sub_wire112(4);
	sub_wire1(16, 5)    <= sub_wire112(5);
	sub_wire1(16, 6)    <= sub_wire112(6);
	sub_wire1(16, 7)    <= sub_wire112(7);
	sub_wire1(16, 8)    <= sub_wire112(8);
	sub_wire1(16, 9)    <= sub_wire112(9);
	sub_wire1(16, 10)    <= sub_wire112(10);
	sub_wire1(16, 11)    <= sub_wire112(11);
	sub_wire1(16, 12)    <= sub_wire112(12);
	sub_wire1(16, 13)    <= sub_wire112(13);
	sub_wire1(16, 14)    <= sub_wire112(14);
	sub_wire1(16, 15)    <= sub_wire112(15);
	sub_wire1(16, 16)    <= sub_wire112(16);
	sub_wire1(16, 17)    <= sub_wire112(17);
	sub_wire1(16, 18)    <= sub_wire112(18);
	sub_wire1(16, 19)    <= sub_wire112(19);
	sub_wire1(16, 20)    <= sub_wire112(20);
	sub_wire1(16, 21)    <= sub_wire112(21);
	sub_wire1(16, 22)    <= sub_wire112(22);
	sub_wire1(16, 23)    <= sub_wire112(23);
	sub_wire1(16, 24)    <= sub_wire112(24);
	sub_wire1(16, 25)    <= sub_wire112(25);
	sub_wire1(16, 26)    <= sub_wire112(26);
	sub_wire1(16, 27)    <= sub_wire112(27);
	sub_wire1(16, 28)    <= sub_wire112(28);
	sub_wire1(16, 29)    <= sub_wire112(29);
	sub_wire1(16, 30)    <= sub_wire112(30);
	sub_wire1(16, 31)    <= sub_wire112(31);
	sub_wire1(15, 0)    <= sub_wire113(0);
	sub_wire1(15, 1)    <= sub_wire113(1);
	sub_wire1(15, 2)    <= sub_wire113(2);
	sub_wire1(15, 3)    <= sub_wire113(3);
	sub_wire1(15, 4)    <= sub_wire113(4);
	sub_wire1(15, 5)    <= sub_wire113(5);
	sub_wire1(15, 6)    <= sub_wire113(6);
	sub_wire1(15, 7)    <= sub_wire113(7);
	sub_wire1(15, 8)    <= sub_wire113(8);
	sub_wire1(15, 9)    <= sub_wire113(9);
	sub_wire1(15, 10)    <= sub_wire113(10);
	sub_wire1(15, 11)    <= sub_wire113(11);
	sub_wire1(15, 12)    <= sub_wire113(12);
	sub_wire1(15, 13)    <= sub_wire113(13);
	sub_wire1(15, 14)    <= sub_wire113(14);
	sub_wire1(15, 15)    <= sub_wire113(15);
	sub_wire1(15, 16)    <= sub_wire113(16);
	sub_wire1(15, 17)    <= sub_wire113(17);
	sub_wire1(15, 18)    <= sub_wire113(18);
	sub_wire1(15, 19)    <= sub_wire113(19);
	sub_wire1(15, 20)    <= sub_wire113(20);
	sub_wire1(15, 21)    <= sub_wire113(21);
	sub_wire1(15, 22)    <= sub_wire113(22);
	sub_wire1(15, 23)    <= sub_wire113(23);
	sub_wire1(15, 24)    <= sub_wire113(24);
	sub_wire1(15, 25)    <= sub_wire113(25);
	sub_wire1(15, 26)    <= sub_wire113(26);
	sub_wire1(15, 27)    <= sub_wire113(27);
	sub_wire1(15, 28)    <= sub_wire113(28);
	sub_wire1(15, 29)    <= sub_wire113(29);
	sub_wire1(15, 30)    <= sub_wire113(30);
	sub_wire1(15, 31)    <= sub_wire113(31);
	sub_wire1(14, 0)    <= sub_wire114(0);
	sub_wire1(14, 1)    <= sub_wire114(1);
	sub_wire1(14, 2)    <= sub_wire114(2);
	sub_wire1(14, 3)    <= sub_wire114(3);
	sub_wire1(14, 4)    <= sub_wire114(4);
	sub_wire1(14, 5)    <= sub_wire114(5);
	sub_wire1(14, 6)    <= sub_wire114(6);
	sub_wire1(14, 7)    <= sub_wire114(7);
	sub_wire1(14, 8)    <= sub_wire114(8);
	sub_wire1(14, 9)    <= sub_wire114(9);
	sub_wire1(14, 10)    <= sub_wire114(10);
	sub_wire1(14, 11)    <= sub_wire114(11);
	sub_wire1(14, 12)    <= sub_wire114(12);
	sub_wire1(14, 13)    <= sub_wire114(13);
	sub_wire1(14, 14)    <= sub_wire114(14);
	sub_wire1(14, 15)    <= sub_wire114(15);
	sub_wire1(14, 16)    <= sub_wire114(16);
	sub_wire1(14, 17)    <= sub_wire114(17);
	sub_wire1(14, 18)    <= sub_wire114(18);
	sub_wire1(14, 19)    <= sub_wire114(19);
	sub_wire1(14, 20)    <= sub_wire114(20);
	sub_wire1(14, 21)    <= sub_wire114(21);
	sub_wire1(14, 22)    <= sub_wire114(22);
	sub_wire1(14, 23)    <= sub_wire114(23);
	sub_wire1(14, 24)    <= sub_wire114(24);
	sub_wire1(14, 25)    <= sub_wire114(25);
	sub_wire1(14, 26)    <= sub_wire114(26);
	sub_wire1(14, 27)    <= sub_wire114(27);
	sub_wire1(14, 28)    <= sub_wire114(28);
	sub_wire1(14, 29)    <= sub_wire114(29);
	sub_wire1(14, 30)    <= sub_wire114(30);
	sub_wire1(14, 31)    <= sub_wire114(31);
	sub_wire1(13, 0)    <= sub_wire115(0);
	sub_wire1(13, 1)    <= sub_wire115(1);
	sub_wire1(13, 2)    <= sub_wire115(2);
	sub_wire1(13, 3)    <= sub_wire115(3);
	sub_wire1(13, 4)    <= sub_wire115(4);
	sub_wire1(13, 5)    <= sub_wire115(5);
	sub_wire1(13, 6)    <= sub_wire115(6);
	sub_wire1(13, 7)    <= sub_wire115(7);
	sub_wire1(13, 8)    <= sub_wire115(8);
	sub_wire1(13, 9)    <= sub_wire115(9);
	sub_wire1(13, 10)    <= sub_wire115(10);
	sub_wire1(13, 11)    <= sub_wire115(11);
	sub_wire1(13, 12)    <= sub_wire115(12);
	sub_wire1(13, 13)    <= sub_wire115(13);
	sub_wire1(13, 14)    <= sub_wire115(14);
	sub_wire1(13, 15)    <= sub_wire115(15);
	sub_wire1(13, 16)    <= sub_wire115(16);
	sub_wire1(13, 17)    <= sub_wire115(17);
	sub_wire1(13, 18)    <= sub_wire115(18);
	sub_wire1(13, 19)    <= sub_wire115(19);
	sub_wire1(13, 20)    <= sub_wire115(20);
	sub_wire1(13, 21)    <= sub_wire115(21);
	sub_wire1(13, 22)    <= sub_wire115(22);
	sub_wire1(13, 23)    <= sub_wire115(23);
	sub_wire1(13, 24)    <= sub_wire115(24);
	sub_wire1(13, 25)    <= sub_wire115(25);
	sub_wire1(13, 26)    <= sub_wire115(26);
	sub_wire1(13, 27)    <= sub_wire115(27);
	sub_wire1(13, 28)    <= sub_wire115(28);
	sub_wire1(13, 29)    <= sub_wire115(29);
	sub_wire1(13, 30)    <= sub_wire115(30);
	sub_wire1(13, 31)    <= sub_wire115(31);
	sub_wire1(12, 0)    <= sub_wire116(0);
	sub_wire1(12, 1)    <= sub_wire116(1);
	sub_wire1(12, 2)    <= sub_wire116(2);
	sub_wire1(12, 3)    <= sub_wire116(3);
	sub_wire1(12, 4)    <= sub_wire116(4);
	sub_wire1(12, 5)    <= sub_wire116(5);
	sub_wire1(12, 6)    <= sub_wire116(6);
	sub_wire1(12, 7)    <= sub_wire116(7);
	sub_wire1(12, 8)    <= sub_wire116(8);
	sub_wire1(12, 9)    <= sub_wire116(9);
	sub_wire1(12, 10)    <= sub_wire116(10);
	sub_wire1(12, 11)    <= sub_wire116(11);
	sub_wire1(12, 12)    <= sub_wire116(12);
	sub_wire1(12, 13)    <= sub_wire116(13);
	sub_wire1(12, 14)    <= sub_wire116(14);
	sub_wire1(12, 15)    <= sub_wire116(15);
	sub_wire1(12, 16)    <= sub_wire116(16);
	sub_wire1(12, 17)    <= sub_wire116(17);
	sub_wire1(12, 18)    <= sub_wire116(18);
	sub_wire1(12, 19)    <= sub_wire116(19);
	sub_wire1(12, 20)    <= sub_wire116(20);
	sub_wire1(12, 21)    <= sub_wire116(21);
	sub_wire1(12, 22)    <= sub_wire116(22);
	sub_wire1(12, 23)    <= sub_wire116(23);
	sub_wire1(12, 24)    <= sub_wire116(24);
	sub_wire1(12, 25)    <= sub_wire116(25);
	sub_wire1(12, 26)    <= sub_wire116(26);
	sub_wire1(12, 27)    <= sub_wire116(27);
	sub_wire1(12, 28)    <= sub_wire116(28);
	sub_wire1(12, 29)    <= sub_wire116(29);
	sub_wire1(12, 30)    <= sub_wire116(30);
	sub_wire1(12, 31)    <= sub_wire116(31);
	sub_wire1(11, 0)    <= sub_wire117(0);
	sub_wire1(11, 1)    <= sub_wire117(1);
	sub_wire1(11, 2)    <= sub_wire117(2);
	sub_wire1(11, 3)    <= sub_wire117(3);
	sub_wire1(11, 4)    <= sub_wire117(4);
	sub_wire1(11, 5)    <= sub_wire117(5);
	sub_wire1(11, 6)    <= sub_wire117(6);
	sub_wire1(11, 7)    <= sub_wire117(7);
	sub_wire1(11, 8)    <= sub_wire117(8);
	sub_wire1(11, 9)    <= sub_wire117(9);
	sub_wire1(11, 10)    <= sub_wire117(10);
	sub_wire1(11, 11)    <= sub_wire117(11);
	sub_wire1(11, 12)    <= sub_wire117(12);
	sub_wire1(11, 13)    <= sub_wire117(13);
	sub_wire1(11, 14)    <= sub_wire117(14);
	sub_wire1(11, 15)    <= sub_wire117(15);
	sub_wire1(11, 16)    <= sub_wire117(16);
	sub_wire1(11, 17)    <= sub_wire117(17);
	sub_wire1(11, 18)    <= sub_wire117(18);
	sub_wire1(11, 19)    <= sub_wire117(19);
	sub_wire1(11, 20)    <= sub_wire117(20);
	sub_wire1(11, 21)    <= sub_wire117(21);
	sub_wire1(11, 22)    <= sub_wire117(22);
	sub_wire1(11, 23)    <= sub_wire117(23);
	sub_wire1(11, 24)    <= sub_wire117(24);
	sub_wire1(11, 25)    <= sub_wire117(25);
	sub_wire1(11, 26)    <= sub_wire117(26);
	sub_wire1(11, 27)    <= sub_wire117(27);
	sub_wire1(11, 28)    <= sub_wire117(28);
	sub_wire1(11, 29)    <= sub_wire117(29);
	sub_wire1(11, 30)    <= sub_wire117(30);
	sub_wire1(11, 31)    <= sub_wire117(31);
	sub_wire1(10, 0)    <= sub_wire118(0);
	sub_wire1(10, 1)    <= sub_wire118(1);
	sub_wire1(10, 2)    <= sub_wire118(2);
	sub_wire1(10, 3)    <= sub_wire118(3);
	sub_wire1(10, 4)    <= sub_wire118(4);
	sub_wire1(10, 5)    <= sub_wire118(5);
	sub_wire1(10, 6)    <= sub_wire118(6);
	sub_wire1(10, 7)    <= sub_wire118(7);
	sub_wire1(10, 8)    <= sub_wire118(8);
	sub_wire1(10, 9)    <= sub_wire118(9);
	sub_wire1(10, 10)    <= sub_wire118(10);
	sub_wire1(10, 11)    <= sub_wire118(11);
	sub_wire1(10, 12)    <= sub_wire118(12);
	sub_wire1(10, 13)    <= sub_wire118(13);
	sub_wire1(10, 14)    <= sub_wire118(14);
	sub_wire1(10, 15)    <= sub_wire118(15);
	sub_wire1(10, 16)    <= sub_wire118(16);
	sub_wire1(10, 17)    <= sub_wire118(17);
	sub_wire1(10, 18)    <= sub_wire118(18);
	sub_wire1(10, 19)    <= sub_wire118(19);
	sub_wire1(10, 20)    <= sub_wire118(20);
	sub_wire1(10, 21)    <= sub_wire118(21);
	sub_wire1(10, 22)    <= sub_wire118(22);
	sub_wire1(10, 23)    <= sub_wire118(23);
	sub_wire1(10, 24)    <= sub_wire118(24);
	sub_wire1(10, 25)    <= sub_wire118(25);
	sub_wire1(10, 26)    <= sub_wire118(26);
	sub_wire1(10, 27)    <= sub_wire118(27);
	sub_wire1(10, 28)    <= sub_wire118(28);
	sub_wire1(10, 29)    <= sub_wire118(29);
	sub_wire1(10, 30)    <= sub_wire118(30);
	sub_wire1(10, 31)    <= sub_wire118(31);
	sub_wire1(9, 0)    <= sub_wire119(0);
	sub_wire1(9, 1)    <= sub_wire119(1);
	sub_wire1(9, 2)    <= sub_wire119(2);
	sub_wire1(9, 3)    <= sub_wire119(3);
	sub_wire1(9, 4)    <= sub_wire119(4);
	sub_wire1(9, 5)    <= sub_wire119(5);
	sub_wire1(9, 6)    <= sub_wire119(6);
	sub_wire1(9, 7)    <= sub_wire119(7);
	sub_wire1(9, 8)    <= sub_wire119(8);
	sub_wire1(9, 9)    <= sub_wire119(9);
	sub_wire1(9, 10)    <= sub_wire119(10);
	sub_wire1(9, 11)    <= sub_wire119(11);
	sub_wire1(9, 12)    <= sub_wire119(12);
	sub_wire1(9, 13)    <= sub_wire119(13);
	sub_wire1(9, 14)    <= sub_wire119(14);
	sub_wire1(9, 15)    <= sub_wire119(15);
	sub_wire1(9, 16)    <= sub_wire119(16);
	sub_wire1(9, 17)    <= sub_wire119(17);
	sub_wire1(9, 18)    <= sub_wire119(18);
	sub_wire1(9, 19)    <= sub_wire119(19);
	sub_wire1(9, 20)    <= sub_wire119(20);
	sub_wire1(9, 21)    <= sub_wire119(21);
	sub_wire1(9, 22)    <= sub_wire119(22);
	sub_wire1(9, 23)    <= sub_wire119(23);
	sub_wire1(9, 24)    <= sub_wire119(24);
	sub_wire1(9, 25)    <= sub_wire119(25);
	sub_wire1(9, 26)    <= sub_wire119(26);
	sub_wire1(9, 27)    <= sub_wire119(27);
	sub_wire1(9, 28)    <= sub_wire119(28);
	sub_wire1(9, 29)    <= sub_wire119(29);
	sub_wire1(9, 30)    <= sub_wire119(30);
	sub_wire1(9, 31)    <= sub_wire119(31);
	sub_wire1(8, 0)    <= sub_wire120(0);
	sub_wire1(8, 1)    <= sub_wire120(1);
	sub_wire1(8, 2)    <= sub_wire120(2);
	sub_wire1(8, 3)    <= sub_wire120(3);
	sub_wire1(8, 4)    <= sub_wire120(4);
	sub_wire1(8, 5)    <= sub_wire120(5);
	sub_wire1(8, 6)    <= sub_wire120(6);
	sub_wire1(8, 7)    <= sub_wire120(7);
	sub_wire1(8, 8)    <= sub_wire120(8);
	sub_wire1(8, 9)    <= sub_wire120(9);
	sub_wire1(8, 10)    <= sub_wire120(10);
	sub_wire1(8, 11)    <= sub_wire120(11);
	sub_wire1(8, 12)    <= sub_wire120(12);
	sub_wire1(8, 13)    <= sub_wire120(13);
	sub_wire1(8, 14)    <= sub_wire120(14);
	sub_wire1(8, 15)    <= sub_wire120(15);
	sub_wire1(8, 16)    <= sub_wire120(16);
	sub_wire1(8, 17)    <= sub_wire120(17);
	sub_wire1(8, 18)    <= sub_wire120(18);
	sub_wire1(8, 19)    <= sub_wire120(19);
	sub_wire1(8, 20)    <= sub_wire120(20);
	sub_wire1(8, 21)    <= sub_wire120(21);
	sub_wire1(8, 22)    <= sub_wire120(22);
	sub_wire1(8, 23)    <= sub_wire120(23);
	sub_wire1(8, 24)    <= sub_wire120(24);
	sub_wire1(8, 25)    <= sub_wire120(25);
	sub_wire1(8, 26)    <= sub_wire120(26);
	sub_wire1(8, 27)    <= sub_wire120(27);
	sub_wire1(8, 28)    <= sub_wire120(28);
	sub_wire1(8, 29)    <= sub_wire120(29);
	sub_wire1(8, 30)    <= sub_wire120(30);
	sub_wire1(8, 31)    <= sub_wire120(31);
	sub_wire1(7, 0)    <= sub_wire121(0);
	sub_wire1(7, 1)    <= sub_wire121(1);
	sub_wire1(7, 2)    <= sub_wire121(2);
	sub_wire1(7, 3)    <= sub_wire121(3);
	sub_wire1(7, 4)    <= sub_wire121(4);
	sub_wire1(7, 5)    <= sub_wire121(5);
	sub_wire1(7, 6)    <= sub_wire121(6);
	sub_wire1(7, 7)    <= sub_wire121(7);
	sub_wire1(7, 8)    <= sub_wire121(8);
	sub_wire1(7, 9)    <= sub_wire121(9);
	sub_wire1(7, 10)    <= sub_wire121(10);
	sub_wire1(7, 11)    <= sub_wire121(11);
	sub_wire1(7, 12)    <= sub_wire121(12);
	sub_wire1(7, 13)    <= sub_wire121(13);
	sub_wire1(7, 14)    <= sub_wire121(14);
	sub_wire1(7, 15)    <= sub_wire121(15);
	sub_wire1(7, 16)    <= sub_wire121(16);
	sub_wire1(7, 17)    <= sub_wire121(17);
	sub_wire1(7, 18)    <= sub_wire121(18);
	sub_wire1(7, 19)    <= sub_wire121(19);
	sub_wire1(7, 20)    <= sub_wire121(20);
	sub_wire1(7, 21)    <= sub_wire121(21);
	sub_wire1(7, 22)    <= sub_wire121(22);
	sub_wire1(7, 23)    <= sub_wire121(23);
	sub_wire1(7, 24)    <= sub_wire121(24);
	sub_wire1(7, 25)    <= sub_wire121(25);
	sub_wire1(7, 26)    <= sub_wire121(26);
	sub_wire1(7, 27)    <= sub_wire121(27);
	sub_wire1(7, 28)    <= sub_wire121(28);
	sub_wire1(7, 29)    <= sub_wire121(29);
	sub_wire1(7, 30)    <= sub_wire121(30);
	sub_wire1(7, 31)    <= sub_wire121(31);
	sub_wire1(6, 0)    <= sub_wire122(0);
	sub_wire1(6, 1)    <= sub_wire122(1);
	sub_wire1(6, 2)    <= sub_wire122(2);
	sub_wire1(6, 3)    <= sub_wire122(3);
	sub_wire1(6, 4)    <= sub_wire122(4);
	sub_wire1(6, 5)    <= sub_wire122(5);
	sub_wire1(6, 6)    <= sub_wire122(6);
	sub_wire1(6, 7)    <= sub_wire122(7);
	sub_wire1(6, 8)    <= sub_wire122(8);
	sub_wire1(6, 9)    <= sub_wire122(9);
	sub_wire1(6, 10)    <= sub_wire122(10);
	sub_wire1(6, 11)    <= sub_wire122(11);
	sub_wire1(6, 12)    <= sub_wire122(12);
	sub_wire1(6, 13)    <= sub_wire122(13);
	sub_wire1(6, 14)    <= sub_wire122(14);
	sub_wire1(6, 15)    <= sub_wire122(15);
	sub_wire1(6, 16)    <= sub_wire122(16);
	sub_wire1(6, 17)    <= sub_wire122(17);
	sub_wire1(6, 18)    <= sub_wire122(18);
	sub_wire1(6, 19)    <= sub_wire122(19);
	sub_wire1(6, 20)    <= sub_wire122(20);
	sub_wire1(6, 21)    <= sub_wire122(21);
	sub_wire1(6, 22)    <= sub_wire122(22);
	sub_wire1(6, 23)    <= sub_wire122(23);
	sub_wire1(6, 24)    <= sub_wire122(24);
	sub_wire1(6, 25)    <= sub_wire122(25);
	sub_wire1(6, 26)    <= sub_wire122(26);
	sub_wire1(6, 27)    <= sub_wire122(27);
	sub_wire1(6, 28)    <= sub_wire122(28);
	sub_wire1(6, 29)    <= sub_wire122(29);
	sub_wire1(6, 30)    <= sub_wire122(30);
	sub_wire1(6, 31)    <= sub_wire122(31);
	sub_wire1(5, 0)    <= sub_wire123(0);
	sub_wire1(5, 1)    <= sub_wire123(1);
	sub_wire1(5, 2)    <= sub_wire123(2);
	sub_wire1(5, 3)    <= sub_wire123(3);
	sub_wire1(5, 4)    <= sub_wire123(4);
	sub_wire1(5, 5)    <= sub_wire123(5);
	sub_wire1(5, 6)    <= sub_wire123(6);
	sub_wire1(5, 7)    <= sub_wire123(7);
	sub_wire1(5, 8)    <= sub_wire123(8);
	sub_wire1(5, 9)    <= sub_wire123(9);
	sub_wire1(5, 10)    <= sub_wire123(10);
	sub_wire1(5, 11)    <= sub_wire123(11);
	sub_wire1(5, 12)    <= sub_wire123(12);
	sub_wire1(5, 13)    <= sub_wire123(13);
	sub_wire1(5, 14)    <= sub_wire123(14);
	sub_wire1(5, 15)    <= sub_wire123(15);
	sub_wire1(5, 16)    <= sub_wire123(16);
	sub_wire1(5, 17)    <= sub_wire123(17);
	sub_wire1(5, 18)    <= sub_wire123(18);
	sub_wire1(5, 19)    <= sub_wire123(19);
	sub_wire1(5, 20)    <= sub_wire123(20);
	sub_wire1(5, 21)    <= sub_wire123(21);
	sub_wire1(5, 22)    <= sub_wire123(22);
	sub_wire1(5, 23)    <= sub_wire123(23);
	sub_wire1(5, 24)    <= sub_wire123(24);
	sub_wire1(5, 25)    <= sub_wire123(25);
	sub_wire1(5, 26)    <= sub_wire123(26);
	sub_wire1(5, 27)    <= sub_wire123(27);
	sub_wire1(5, 28)    <= sub_wire123(28);
	sub_wire1(5, 29)    <= sub_wire123(29);
	sub_wire1(5, 30)    <= sub_wire123(30);
	sub_wire1(5, 31)    <= sub_wire123(31);
	sub_wire1(4, 0)    <= sub_wire124(0);
	sub_wire1(4, 1)    <= sub_wire124(1);
	sub_wire1(4, 2)    <= sub_wire124(2);
	sub_wire1(4, 3)    <= sub_wire124(3);
	sub_wire1(4, 4)    <= sub_wire124(4);
	sub_wire1(4, 5)    <= sub_wire124(5);
	sub_wire1(4, 6)    <= sub_wire124(6);
	sub_wire1(4, 7)    <= sub_wire124(7);
	sub_wire1(4, 8)    <= sub_wire124(8);
	sub_wire1(4, 9)    <= sub_wire124(9);
	sub_wire1(4, 10)    <= sub_wire124(10);
	sub_wire1(4, 11)    <= sub_wire124(11);
	sub_wire1(4, 12)    <= sub_wire124(12);
	sub_wire1(4, 13)    <= sub_wire124(13);
	sub_wire1(4, 14)    <= sub_wire124(14);
	sub_wire1(4, 15)    <= sub_wire124(15);
	sub_wire1(4, 16)    <= sub_wire124(16);
	sub_wire1(4, 17)    <= sub_wire124(17);
	sub_wire1(4, 18)    <= sub_wire124(18);
	sub_wire1(4, 19)    <= sub_wire124(19);
	sub_wire1(4, 20)    <= sub_wire124(20);
	sub_wire1(4, 21)    <= sub_wire124(21);
	sub_wire1(4, 22)    <= sub_wire124(22);
	sub_wire1(4, 23)    <= sub_wire124(23);
	sub_wire1(4, 24)    <= sub_wire124(24);
	sub_wire1(4, 25)    <= sub_wire124(25);
	sub_wire1(4, 26)    <= sub_wire124(26);
	sub_wire1(4, 27)    <= sub_wire124(27);
	sub_wire1(4, 28)    <= sub_wire124(28);
	sub_wire1(4, 29)    <= sub_wire124(29);
	sub_wire1(4, 30)    <= sub_wire124(30);
	sub_wire1(4, 31)    <= sub_wire124(31);
	sub_wire1(3, 0)    <= sub_wire125(0);
	sub_wire1(3, 1)    <= sub_wire125(1);
	sub_wire1(3, 2)    <= sub_wire125(2);
	sub_wire1(3, 3)    <= sub_wire125(3);
	sub_wire1(3, 4)    <= sub_wire125(4);
	sub_wire1(3, 5)    <= sub_wire125(5);
	sub_wire1(3, 6)    <= sub_wire125(6);
	sub_wire1(3, 7)    <= sub_wire125(7);
	sub_wire1(3, 8)    <= sub_wire125(8);
	sub_wire1(3, 9)    <= sub_wire125(9);
	sub_wire1(3, 10)    <= sub_wire125(10);
	sub_wire1(3, 11)    <= sub_wire125(11);
	sub_wire1(3, 12)    <= sub_wire125(12);
	sub_wire1(3, 13)    <= sub_wire125(13);
	sub_wire1(3, 14)    <= sub_wire125(14);
	sub_wire1(3, 15)    <= sub_wire125(15);
	sub_wire1(3, 16)    <= sub_wire125(16);
	sub_wire1(3, 17)    <= sub_wire125(17);
	sub_wire1(3, 18)    <= sub_wire125(18);
	sub_wire1(3, 19)    <= sub_wire125(19);
	sub_wire1(3, 20)    <= sub_wire125(20);
	sub_wire1(3, 21)    <= sub_wire125(21);
	sub_wire1(3, 22)    <= sub_wire125(22);
	sub_wire1(3, 23)    <= sub_wire125(23);
	sub_wire1(3, 24)    <= sub_wire125(24);
	sub_wire1(3, 25)    <= sub_wire125(25);
	sub_wire1(3, 26)    <= sub_wire125(26);
	sub_wire1(3, 27)    <= sub_wire125(27);
	sub_wire1(3, 28)    <= sub_wire125(28);
	sub_wire1(3, 29)    <= sub_wire125(29);
	sub_wire1(3, 30)    <= sub_wire125(30);
	sub_wire1(3, 31)    <= sub_wire125(31);
	sub_wire1(2, 0)    <= sub_wire126(0);
	sub_wire1(2, 1)    <= sub_wire126(1);
	sub_wire1(2, 2)    <= sub_wire126(2);
	sub_wire1(2, 3)    <= sub_wire126(3);
	sub_wire1(2, 4)    <= sub_wire126(4);
	sub_wire1(2, 5)    <= sub_wire126(5);
	sub_wire1(2, 6)    <= sub_wire126(6);
	sub_wire1(2, 7)    <= sub_wire126(7);
	sub_wire1(2, 8)    <= sub_wire126(8);
	sub_wire1(2, 9)    <= sub_wire126(9);
	sub_wire1(2, 10)    <= sub_wire126(10);
	sub_wire1(2, 11)    <= sub_wire126(11);
	sub_wire1(2, 12)    <= sub_wire126(12);
	sub_wire1(2, 13)    <= sub_wire126(13);
	sub_wire1(2, 14)    <= sub_wire126(14);
	sub_wire1(2, 15)    <= sub_wire126(15);
	sub_wire1(2, 16)    <= sub_wire126(16);
	sub_wire1(2, 17)    <= sub_wire126(17);
	sub_wire1(2, 18)    <= sub_wire126(18);
	sub_wire1(2, 19)    <= sub_wire126(19);
	sub_wire1(2, 20)    <= sub_wire126(20);
	sub_wire1(2, 21)    <= sub_wire126(21);
	sub_wire1(2, 22)    <= sub_wire126(22);
	sub_wire1(2, 23)    <= sub_wire126(23);
	sub_wire1(2, 24)    <= sub_wire126(24);
	sub_wire1(2, 25)    <= sub_wire126(25);
	sub_wire1(2, 26)    <= sub_wire126(26);
	sub_wire1(2, 27)    <= sub_wire126(27);
	sub_wire1(2, 28)    <= sub_wire126(28);
	sub_wire1(2, 29)    <= sub_wire126(29);
	sub_wire1(2, 30)    <= sub_wire126(30);
	sub_wire1(2, 31)    <= sub_wire126(31);
	sub_wire1(1, 0)    <= sub_wire127(0);
	sub_wire1(1, 1)    <= sub_wire127(1);
	sub_wire1(1, 2)    <= sub_wire127(2);
	sub_wire1(1, 3)    <= sub_wire127(3);
	sub_wire1(1, 4)    <= sub_wire127(4);
	sub_wire1(1, 5)    <= sub_wire127(5);
	sub_wire1(1, 6)    <= sub_wire127(6);
	sub_wire1(1, 7)    <= sub_wire127(7);
	sub_wire1(1, 8)    <= sub_wire127(8);
	sub_wire1(1, 9)    <= sub_wire127(9);
	sub_wire1(1, 10)    <= sub_wire127(10);
	sub_wire1(1, 11)    <= sub_wire127(11);
	sub_wire1(1, 12)    <= sub_wire127(12);
	sub_wire1(1, 13)    <= sub_wire127(13);
	sub_wire1(1, 14)    <= sub_wire127(14);
	sub_wire1(1, 15)    <= sub_wire127(15);
	sub_wire1(1, 16)    <= sub_wire127(16);
	sub_wire1(1, 17)    <= sub_wire127(17);
	sub_wire1(1, 18)    <= sub_wire127(18);
	sub_wire1(1, 19)    <= sub_wire127(19);
	sub_wire1(1, 20)    <= sub_wire127(20);
	sub_wire1(1, 21)    <= sub_wire127(21);
	sub_wire1(1, 22)    <= sub_wire127(22);
	sub_wire1(1, 23)    <= sub_wire127(23);
	sub_wire1(1, 24)    <= sub_wire127(24);
	sub_wire1(1, 25)    <= sub_wire127(25);
	sub_wire1(1, 26)    <= sub_wire127(26);
	sub_wire1(1, 27)    <= sub_wire127(27);
	sub_wire1(1, 28)    <= sub_wire127(28);
	sub_wire1(1, 29)    <= sub_wire127(29);
	sub_wire1(1, 30)    <= sub_wire127(30);
	sub_wire1(1, 31)    <= sub_wire127(31);
	sub_wire1(0, 0)    <= sub_wire128(0);
	sub_wire1(0, 1)    <= sub_wire128(1);
	sub_wire1(0, 2)    <= sub_wire128(2);
	sub_wire1(0, 3)    <= sub_wire128(3);
	sub_wire1(0, 4)    <= sub_wire128(4);
	sub_wire1(0, 5)    <= sub_wire128(5);
	sub_wire1(0, 6)    <= sub_wire128(6);
	sub_wire1(0, 7)    <= sub_wire128(7);
	sub_wire1(0, 8)    <= sub_wire128(8);
	sub_wire1(0, 9)    <= sub_wire128(9);
	sub_wire1(0, 10)    <= sub_wire128(10);
	sub_wire1(0, 11)    <= sub_wire128(11);
	sub_wire1(0, 12)    <= sub_wire128(12);
	sub_wire1(0, 13)    <= sub_wire128(13);
	sub_wire1(0, 14)    <= sub_wire128(14);
	sub_wire1(0, 15)    <= sub_wire128(15);
	sub_wire1(0, 16)    <= sub_wire128(16);
	sub_wire1(0, 17)    <= sub_wire128(17);
	sub_wire1(0, 18)    <= sub_wire128(18);
	sub_wire1(0, 19)    <= sub_wire128(19);
	sub_wire1(0, 20)    <= sub_wire128(20);
	sub_wire1(0, 21)    <= sub_wire128(21);
	sub_wire1(0, 22)    <= sub_wire128(22);
	sub_wire1(0, 23)    <= sub_wire128(23);
	sub_wire1(0, 24)    <= sub_wire128(24);
	sub_wire1(0, 25)    <= sub_wire128(25);
	sub_wire1(0, 26)    <= sub_wire128(26);
	sub_wire1(0, 27)    <= sub_wire128(27);
	sub_wire1(0, 28)    <= sub_wire128(28);
	sub_wire1(0, 29)    <= sub_wire128(29);
	sub_wire1(0, 30)    <= sub_wire128(30);
	sub_wire1(0, 31)    <= sub_wire128(31);
	result    <= sub_wire129(31 DOWNTO 0);

	LPM_MUX_component : LPM_MUX
	GENERIC MAP (
		lpm_size => 128,
		lpm_type => "LPM_MUX",
		lpm_width => 32,
		lpm_widths => 7
	)
	PORT MAP (
		data => sub_wire1,
		sel => sel,
		result => sub_wire129
	);



END SYN;

-- ============================================================
-- CNX file retrieval info
-- ============================================================
-- Retrieval info: PRIVATE: INTENDED_DEVICE_FAMILY STRING "Cyclone IV E"
-- Retrieval info: PRIVATE: SYNTH_WRAPPER_GEN_POSTFIX STRING "0"
-- Retrieval info: PRIVATE: new_diagram STRING "1"
-- Retrieval info: LIBRARY: lpm lpm.lpm_components.all
-- Retrieval info: CONSTANT: LPM_SIZE NUMERIC "128"
-- Retrieval info: CONSTANT: LPM_TYPE STRING "LPM_MUX"
-- Retrieval info: CONSTANT: LPM_WIDTH NUMERIC "32"
-- Retrieval info: CONSTANT: LPM_WIDTHS NUMERIC "7"
-- Retrieval info: USED_PORT: data0x 0 0 32 0 INPUT NODEFVAL "data0x[31..0]"
-- Retrieval info: USED_PORT: data100x 0 0 32 0 INPUT NODEFVAL "data100x[31..0]"
-- Retrieval info: USED_PORT: data101x 0 0 32 0 INPUT NODEFVAL "data101x[31..0]"
-- Retrieval info: USED_PORT: data102x 0 0 32 0 INPUT NODEFVAL "data102x[31..0]"
-- Retrieval info: USED_PORT: data103x 0 0 32 0 INPUT NODEFVAL "data103x[31..0]"
-- Retrieval info: USED_PORT: data104x 0 0 32 0 INPUT NODEFVAL "data104x[31..0]"
-- Retrieval info: USED_PORT: data105x 0 0 32 0 INPUT NODEFVAL "data105x[31..0]"
-- Retrieval info: USED_PORT: data106x 0 0 32 0 INPUT NODEFVAL "data106x[31..0]"
-- Retrieval info: USED_PORT: data107x 0 0 32 0 INPUT NODEFVAL "data107x[31..0]"
-- Retrieval info: USED_PORT: data108x 0 0 32 0 INPUT NODEFVAL "data108x[31..0]"
-- Retrieval info: USED_PORT: data109x 0 0 32 0 INPUT NODEFVAL "data109x[31..0]"
-- Retrieval info: USED_PORT: data10x 0 0 32 0 INPUT NODEFVAL "data10x[31..0]"
-- Retrieval info: USED_PORT: data110x 0 0 32 0 INPUT NODEFVAL "data110x[31..0]"
-- Retrieval info: USED_PORT: data111x 0 0 32 0 INPUT NODEFVAL "data111x[31..0]"
-- Retrieval info: USED_PORT: data112x 0 0 32 0 INPUT NODEFVAL "data112x[31..0]"
-- Retrieval info: USED_PORT: data113x 0 0 32 0 INPUT NODEFVAL "data113x[31..0]"
-- Retrieval info: USED_PORT: data114x 0 0 32 0 INPUT NODEFVAL "data114x[31..0]"
-- Retrieval info: USED_PORT: data115x 0 0 32 0 INPUT NODEFVAL "data115x[31..0]"
-- Retrieval info: USED_PORT: data116x 0 0 32 0 INPUT NODEFVAL "data116x[31..0]"
-- Retrieval info: USED_PORT: data117x 0 0 32 0 INPUT NODEFVAL "data117x[31..0]"
-- Retrieval info: USED_PORT: data118x 0 0 32 0 INPUT NODEFVAL "data118x[31..0]"
-- Retrieval info: USED_PORT: data119x 0 0 32 0 INPUT NODEFVAL "data119x[31..0]"
-- Retrieval info: USED_PORT: data11x 0 0 32 0 INPUT NODEFVAL "data11x[31..0]"
-- Retrieval info: USED_PORT: data120x 0 0 32 0 INPUT NODEFVAL "data120x[31..0]"
-- Retrieval info: USED_PORT: data121x 0 0 32 0 INPUT NODEFVAL "data121x[31..0]"
-- Retrieval info: USED_PORT: data122x 0 0 32 0 INPUT NODEFVAL "data122x[31..0]"
-- Retrieval info: USED_PORT: data123x 0 0 32 0 INPUT NODEFVAL "data123x[31..0]"
-- Retrieval info: USED_PORT: data124x 0 0 32 0 INPUT NODEFVAL "data124x[31..0]"
-- Retrieval info: USED_PORT: data125x 0 0 32 0 INPUT NODEFVAL "data125x[31..0]"
-- Retrieval info: USED_PORT: data126x 0 0 32 0 INPUT NODEFVAL "data126x[31..0]"
-- Retrieval info: USED_PORT: data127x 0 0 32 0 INPUT NODEFVAL "data127x[31..0]"
-- Retrieval info: USED_PORT: data12x 0 0 32 0 INPUT NODEFVAL "data12x[31..0]"
-- Retrieval info: USED_PORT: data13x 0 0 32 0 INPUT NODEFVAL "data13x[31..0]"
-- Retrieval info: USED_PORT: data14x 0 0 32 0 INPUT NODEFVAL "data14x[31..0]"
-- Retrieval info: USED_PORT: data15x 0 0 32 0 INPUT NODEFVAL "data15x[31..0]"
-- Retrieval info: USED_PORT: data16x 0 0 32 0 INPUT NODEFVAL "data16x[31..0]"
-- Retrieval info: USED_PORT: data17x 0 0 32 0 INPUT NODEFVAL "data17x[31..0]"
-- Retrieval info: USED_PORT: data18x 0 0 32 0 INPUT NODEFVAL "data18x[31..0]"
-- Retrieval info: USED_PORT: data19x 0 0 32 0 INPUT NODEFVAL "data19x[31..0]"
-- Retrieval info: USED_PORT: data1x 0 0 32 0 INPUT NODEFVAL "data1x[31..0]"
-- Retrieval info: USED_PORT: data20x 0 0 32 0 INPUT NODEFVAL "data20x[31..0]"
-- Retrieval info: USED_PORT: data21x 0 0 32 0 INPUT NODEFVAL "data21x[31..0]"
-- Retrieval info: USED_PORT: data22x 0 0 32 0 INPUT NODEFVAL "data22x[31..0]"
-- Retrieval info: USED_PORT: data23x 0 0 32 0 INPUT NODEFVAL "data23x[31..0]"
-- Retrieval info: USED_PORT: data24x 0 0 32 0 INPUT NODEFVAL "data24x[31..0]"
-- Retrieval info: USED_PORT: data25x 0 0 32 0 INPUT NODEFVAL "data25x[31..0]"
-- Retrieval info: USED_PORT: data26x 0 0 32 0 INPUT NODEFVAL "data26x[31..0]"
-- Retrieval info: USED_PORT: data27x 0 0 32 0 INPUT NODEFVAL "data27x[31..0]"
-- Retrieval info: USED_PORT: data28x 0 0 32 0 INPUT NODEFVAL "data28x[31..0]"
-- Retrieval info: USED_PORT: data29x 0 0 32 0 INPUT NODEFVAL "data29x[31..0]"
-- Retrieval info: USED_PORT: data2x 0 0 32 0 INPUT NODEFVAL "data2x[31..0]"
-- Retrieval info: USED_PORT: data30x 0 0 32 0 INPUT NODEFVAL "data30x[31..0]"
-- Retrieval info: USED_PORT: data31x 0 0 32 0 INPUT NODEFVAL "data31x[31..0]"
-- Retrieval info: USED_PORT: data32x 0 0 32 0 INPUT NODEFVAL "data32x[31..0]"
-- Retrieval info: USED_PORT: data33x 0 0 32 0 INPUT NODEFVAL "data33x[31..0]"
-- Retrieval info: USED_PORT: data34x 0 0 32 0 INPUT NODEFVAL "data34x[31..0]"
-- Retrieval info: USED_PORT: data35x 0 0 32 0 INPUT NODEFVAL "data35x[31..0]"
-- Retrieval info: USED_PORT: data36x 0 0 32 0 INPUT NODEFVAL "data36x[31..0]"
-- Retrieval info: USED_PORT: data37x 0 0 32 0 INPUT NODEFVAL "data37x[31..0]"
-- Retrieval info: USED_PORT: data38x 0 0 32 0 INPUT NODEFVAL "data38x[31..0]"
-- Retrieval info: USED_PORT: data39x 0 0 32 0 INPUT NODEFVAL "data39x[31..0]"
-- Retrieval info: USED_PORT: data3x 0 0 32 0 INPUT NODEFVAL "data3x[31..0]"
-- Retrieval info: USED_PORT: data40x 0 0 32 0 INPUT NODEFVAL "data40x[31..0]"
-- Retrieval info: USED_PORT: data41x 0 0 32 0 INPUT NODEFVAL "data41x[31..0]"
-- Retrieval info: USED_PORT: data42x 0 0 32 0 INPUT NODEFVAL "data42x[31..0]"
-- Retrieval info: USED_PORT: data43x 0 0 32 0 INPUT NODEFVAL "data43x[31..0]"
-- Retrieval info: USED_PORT: data44x 0 0 32 0 INPUT NODEFVAL "data44x[31..0]"
-- Retrieval info: USED_PORT: data45x 0 0 32 0 INPUT NODEFVAL "data45x[31..0]"
-- Retrieval info: USED_PORT: data46x 0 0 32 0 INPUT NODEFVAL "data46x[31..0]"
-- Retrieval info: USED_PORT: data47x 0 0 32 0 INPUT NODEFVAL "data47x[31..0]"
-- Retrieval info: USED_PORT: data48x 0 0 32 0 INPUT NODEFVAL "data48x[31..0]"
-- Retrieval info: USED_PORT: data49x 0 0 32 0 INPUT NODEFVAL "data49x[31..0]"
-- Retrieval info: USED_PORT: data4x 0 0 32 0 INPUT NODEFVAL "data4x[31..0]"
-- Retrieval info: USED_PORT: data50x 0 0 32 0 INPUT NODEFVAL "data50x[31..0]"
-- Retrieval info: USED_PORT: data51x 0 0 32 0 INPUT NODEFVAL "data51x[31..0]"
-- Retrieval info: USED_PORT: data52x 0 0 32 0 INPUT NODEFVAL "data52x[31..0]"
-- Retrieval info: USED_PORT: data53x 0 0 32 0 INPUT NODEFVAL "data53x[31..0]"
-- Retrieval info: USED_PORT: data54x 0 0 32 0 INPUT NODEFVAL "data54x[31..0]"
-- Retrieval info: USED_PORT: data55x 0 0 32 0 INPUT NODEFVAL "data55x[31..0]"
-- Retrieval info: USED_PORT: data56x 0 0 32 0 INPUT NODEFVAL "data56x[31..0]"
-- Retrieval info: USED_PORT: data57x 0 0 32 0 INPUT NODEFVAL "data57x[31..0]"
-- Retrieval info: USED_PORT: data58x 0 0 32 0 INPUT NODEFVAL "data58x[31..0]"
-- Retrieval info: USED_PORT: data59x 0 0 32 0 INPUT NODEFVAL "data59x[31..0]"
-- Retrieval info: USED_PORT: data5x 0 0 32 0 INPUT NODEFVAL "data5x[31..0]"
-- Retrieval info: USED_PORT: data60x 0 0 32 0 INPUT NODEFVAL "data60x[31..0]"
-- Retrieval info: USED_PORT: data61x 0 0 32 0 INPUT NODEFVAL "data61x[31..0]"
-- Retrieval info: USED_PORT: data62x 0 0 32 0 INPUT NODEFVAL "data62x[31..0]"
-- Retrieval info: USED_PORT: data63x 0 0 32 0 INPUT NODEFVAL "data63x[31..0]"
-- Retrieval info: USED_PORT: data64x 0 0 32 0 INPUT NODEFVAL "data64x[31..0]"
-- Retrieval info: USED_PORT: data65x 0 0 32 0 INPUT NODEFVAL "data65x[31..0]"
-- Retrieval info: USED_PORT: data66x 0 0 32 0 INPUT NODEFVAL "data66x[31..0]"
-- Retrieval info: USED_PORT: data67x 0 0 32 0 INPUT NODEFVAL "data67x[31..0]"
-- Retrieval info: USED_PORT: data68x 0 0 32 0 INPUT NODEFVAL "data68x[31..0]"
-- Retrieval info: USED_PORT: data69x 0 0 32 0 INPUT NODEFVAL "data69x[31..0]"
-- Retrieval info: USED_PORT: data6x 0 0 32 0 INPUT NODEFVAL "data6x[31..0]"
-- Retrieval info: USED_PORT: data70x 0 0 32 0 INPUT NODEFVAL "data70x[31..0]"
-- Retrieval info: USED_PORT: data71x 0 0 32 0 INPUT NODEFVAL "data71x[31..0]"
-- Retrieval info: USED_PORT: data72x 0 0 32 0 INPUT NODEFVAL "data72x[31..0]"
-- Retrieval info: USED_PORT: data73x 0 0 32 0 INPUT NODEFVAL "data73x[31..0]"
-- Retrieval info: USED_PORT: data74x 0 0 32 0 INPUT NODEFVAL "data74x[31..0]"
-- Retrieval info: USED_PORT: data75x 0 0 32 0 INPUT NODEFVAL "data75x[31..0]"
-- Retrieval info: USED_PORT: data76x 0 0 32 0 INPUT NODEFVAL "data76x[31..0]"
-- Retrieval info: USED_PORT: data77x 0 0 32 0 INPUT NODEFVAL "data77x[31..0]"
-- Retrieval info: USED_PORT: data78x 0 0 32 0 INPUT NODEFVAL "data78x[31..0]"
-- Retrieval info: USED_PORT: data79x 0 0 32 0 INPUT NODEFVAL "data79x[31..0]"
-- Retrieval info: USED_PORT: data7x 0 0 32 0 INPUT NODEFVAL "data7x[31..0]"
-- Retrieval info: USED_PORT: data80x 0 0 32 0 INPUT NODEFVAL "data80x[31..0]"
-- Retrieval info: USED_PORT: data81x 0 0 32 0 INPUT NODEFVAL "data81x[31..0]"
-- Retrieval info: USED_PORT: data82x 0 0 32 0 INPUT NODEFVAL "data82x[31..0]"
-- Retrieval info: USED_PORT: data83x 0 0 32 0 INPUT NODEFVAL "data83x[31..0]"
-- Retrieval info: USED_PORT: data84x 0 0 32 0 INPUT NODEFVAL "data84x[31..0]"
-- Retrieval info: USED_PORT: data85x 0 0 32 0 INPUT NODEFVAL "data85x[31..0]"
-- Retrieval info: USED_PORT: data86x 0 0 32 0 INPUT NODEFVAL "data86x[31..0]"
-- Retrieval info: USED_PORT: data87x 0 0 32 0 INPUT NODEFVAL "data87x[31..0]"
-- Retrieval info: USED_PORT: data88x 0 0 32 0 INPUT NODEFVAL "data88x[31..0]"
-- Retrieval info: USED_PORT: data89x 0 0 32 0 INPUT NODEFVAL "data89x[31..0]"
-- Retrieval info: USED_PORT: data8x 0 0 32 0 INPUT NODEFVAL "data8x[31..0]"
-- Retrieval info: USED_PORT: data90x 0 0 32 0 INPUT NODEFVAL "data90x[31..0]"
-- Retrieval info: USED_PORT: data91x 0 0 32 0 INPUT NODEFVAL "data91x[31..0]"
-- Retrieval info: USED_PORT: data92x 0 0 32 0 INPUT NODEFVAL "data92x[31..0]"
-- Retrieval info: USED_PORT: data93x 0 0 32 0 INPUT NODEFVAL "data93x[31..0]"
-- Retrieval info: USED_PORT: data94x 0 0 32 0 INPUT NODEFVAL "data94x[31..0]"
-- Retrieval info: USED_PORT: data95x 0 0 32 0 INPUT NODEFVAL "data95x[31..0]"
-- Retrieval info: USED_PORT: data96x 0 0 32 0 INPUT NODEFVAL "data96x[31..0]"
-- Retrieval info: USED_PORT: data97x 0 0 32 0 INPUT NODEFVAL "data97x[31..0]"
-- Retrieval info: USED_PORT: data98x 0 0 32 0 INPUT NODEFVAL "data98x[31..0]"
-- Retrieval info: USED_PORT: data99x 0 0 32 0 INPUT NODEFVAL "data99x[31..0]"
-- Retrieval info: USED_PORT: data9x 0 0 32 0 INPUT NODEFVAL "data9x[31..0]"
-- Retrieval info: USED_PORT: result 0 0 32 0 OUTPUT NODEFVAL "result[31..0]"
-- Retrieval info: USED_PORT: sel 0 0 7 0 INPUT NODEFVAL "sel[6..0]"
-- Retrieval info: CONNECT: @data 1 0 32 0 data0x 0 0 32 0
-- Retrieval info: CONNECT: @data 1 100 32 0 data100x 0 0 32 0
-- Retrieval info: CONNECT: @data 1 101 32 0 data101x 0 0 32 0
-- Retrieval info: CONNECT: @data 1 102 32 0 data102x 0 0 32 0
-- Retrieval info: CONNECT: @data 1 103 32 0 data103x 0 0 32 0
-- Retrieval info: CONNECT: @data 1 104 32 0 data104x 0 0 32 0
-- Retrieval info: CONNECT: @data 1 105 32 0 data105x 0 0 32 0
-- Retrieval info: CONNECT: @data 1 106 32 0 data106x 0 0 32 0
-- Retrieval info: CONNECT: @data 1 107 32 0 data107x 0 0 32 0
-- Retrieval info: CONNECT: @data 1 108 32 0 data108x 0 0 32 0
-- Retrieval info: CONNECT: @data 1 109 32 0 data109x 0 0 32 0
-- Retrieval info: CONNECT: @data 1 10 32 0 data10x 0 0 32 0
-- Retrieval info: CONNECT: @data 1 110 32 0 data110x 0 0 32 0
-- Retrieval info: CONNECT: @data 1 111 32 0 data111x 0 0 32 0
-- Retrieval info: CONNECT: @data 1 112 32 0 data112x 0 0 32 0
-- Retrieval info: CONNECT: @data 1 113 32 0 data113x 0 0 32 0
-- Retrieval info: CONNECT: @data 1 114 32 0 data114x 0 0 32 0
-- Retrieval info: CONNECT: @data 1 115 32 0 data115x 0 0 32 0
-- Retrieval info: CONNECT: @data 1 116 32 0 data116x 0 0 32 0
-- Retrieval info: CONNECT: @data 1 117 32 0 data117x 0 0 32 0
-- Retrieval info: CONNECT: @data 1 118 32 0 data118x 0 0 32 0
-- Retrieval info: CONNECT: @data 1 119 32 0 data119x 0 0 32 0
-- Retrieval info: CONNECT: @data 1 11 32 0 data11x 0 0 32 0
-- Retrieval info: CONNECT: @data 1 120 32 0 data120x 0 0 32 0
-- Retrieval info: CONNECT: @data 1 121 32 0 data121x 0 0 32 0
-- Retrieval info: CONNECT: @data 1 122 32 0 data122x 0 0 32 0
-- Retrieval info: CONNECT: @data 1 123 32 0 data123x 0 0 32 0
-- Retrieval info: CONNECT: @data 1 124 32 0 data124x 0 0 32 0
-- Retrieval info: CONNECT: @data 1 125 32 0 data125x 0 0 32 0
-- Retrieval info: CONNECT: @data 1 126 32 0 data126x 0 0 32 0
-- Retrieval info: CONNECT: @data 1 127 32 0 data127x 0 0 32 0
-- Retrieval info: CONNECT: @data 1 12 32 0 data12x 0 0 32 0
-- Retrieval info: CONNECT: @data 1 13 32 0 data13x 0 0 32 0
-- Retrieval info: CONNECT: @data 1 14 32 0 data14x 0 0 32 0
-- Retrieval info: CONNECT: @data 1 15 32 0 data15x 0 0 32 0
-- Retrieval info: CONNECT: @data 1 16 32 0 data16x 0 0 32 0
-- Retrieval info: CONNECT: @data 1 17 32 0 data17x 0 0 32 0
-- Retrieval info: CONNECT: @data 1 18 32 0 data18x 0 0 32 0
-- Retrieval info: CONNECT: @data 1 19 32 0 data19x 0 0 32 0
-- Retrieval info: CONNECT: @data 1 1 32 0 data1x 0 0 32 0
-- Retrieval info: CONNECT: @data 1 20 32 0 data20x 0 0 32 0
-- Retrieval info: CONNECT: @data 1 21 32 0 data21x 0 0 32 0
-- Retrieval info: CONNECT: @data 1 22 32 0 data22x 0 0 32 0
-- Retrieval info: CONNECT: @data 1 23 32 0 data23x 0 0 32 0
-- Retrieval info: CONNECT: @data 1 24 32 0 data24x 0 0 32 0
-- Retrieval info: CONNECT: @data 1 25 32 0 data25x 0 0 32 0
-- Retrieval info: CONNECT: @data 1 26 32 0 data26x 0 0 32 0
-- Retrieval info: CONNECT: @data 1 27 32 0 data27x 0 0 32 0
-- Retrieval info: CONNECT: @data 1 28 32 0 data28x 0 0 32 0
-- Retrieval info: CONNECT: @data 1 29 32 0 data29x 0 0 32 0
-- Retrieval info: CONNECT: @data 1 2 32 0 data2x 0 0 32 0
-- Retrieval info: CONNECT: @data 1 30 32 0 data30x 0 0 32 0
-- Retrieval info: CONNECT: @data 1 31 32 0 data31x 0 0 32 0
-- Retrieval info: CONNECT: @data 1 32 32 0 data32x 0 0 32 0
-- Retrieval info: CONNECT: @data 1 33 32 0 data33x 0 0 32 0
-- Retrieval info: CONNECT: @data 1 34 32 0 data34x 0 0 32 0
-- Retrieval info: CONNECT: @data 1 35 32 0 data35x 0 0 32 0
-- Retrieval info: CONNECT: @data 1 36 32 0 data36x 0 0 32 0
-- Retrieval info: CONNECT: @data 1 37 32 0 data37x 0 0 32 0
-- Retrieval info: CONNECT: @data 1 38 32 0 data38x 0 0 32 0
-- Retrieval info: CONNECT: @data 1 39 32 0 data39x 0 0 32 0
-- Retrieval info: CONNECT: @data 1 3 32 0 data3x 0 0 32 0
-- Retrieval info: CONNECT: @data 1 40 32 0 data40x 0 0 32 0
-- Retrieval info: CONNECT: @data 1 41 32 0 data41x 0 0 32 0
-- Retrieval info: CONNECT: @data 1 42 32 0 data42x 0 0 32 0
-- Retrieval info: CONNECT: @data 1 43 32 0 data43x 0 0 32 0
-- Retrieval info: CONNECT: @data 1 44 32 0 data44x 0 0 32 0
-- Retrieval info: CONNECT: @data 1 45 32 0 data45x 0 0 32 0
-- Retrieval info: CONNECT: @data 1 46 32 0 data46x 0 0 32 0
-- Retrieval info: CONNECT: @data 1 47 32 0 data47x 0 0 32 0
-- Retrieval info: CONNECT: @data 1 48 32 0 data48x 0 0 32 0
-- Retrieval info: CONNECT: @data 1 49 32 0 data49x 0 0 32 0
-- Retrieval info: CONNECT: @data 1 4 32 0 data4x 0 0 32 0
-- Retrieval info: CONNECT: @data 1 50 32 0 data50x 0 0 32 0
-- Retrieval info: CONNECT: @data 1 51 32 0 data51x 0 0 32 0
-- Retrieval info: CONNECT: @data 1 52 32 0 data52x 0 0 32 0
-- Retrieval info: CONNECT: @data 1 53 32 0 data53x 0 0 32 0
-- Retrieval info: CONNECT: @data 1 54 32 0 data54x 0 0 32 0
-- Retrieval info: CONNECT: @data 1 55 32 0 data55x 0 0 32 0
-- Retrieval info: CONNECT: @data 1 56 32 0 data56x 0 0 32 0
-- Retrieval info: CONNECT: @data 1 57 32 0 data57x 0 0 32 0
-- Retrieval info: CONNECT: @data 1 58 32 0 data58x 0 0 32 0
-- Retrieval info: CONNECT: @data 1 59 32 0 data59x 0 0 32 0
-- Retrieval info: CONNECT: @data 1 5 32 0 data5x 0 0 32 0
-- Retrieval info: CONNECT: @data 1 60 32 0 data60x 0 0 32 0
-- Retrieval info: CONNECT: @data 1 61 32 0 data61x 0 0 32 0
-- Retrieval info: CONNECT: @data 1 62 32 0 data62x 0 0 32 0
-- Retrieval info: CONNECT: @data 1 63 32 0 data63x 0 0 32 0
-- Retrieval info: CONNECT: @data 1 64 32 0 data64x 0 0 32 0
-- Retrieval info: CONNECT: @data 1 65 32 0 data65x 0 0 32 0
-- Retrieval info: CONNECT: @data 1 66 32 0 data66x 0 0 32 0
-- Retrieval info: CONNECT: @data 1 67 32 0 data67x 0 0 32 0
-- Retrieval info: CONNECT: @data 1 68 32 0 data68x 0 0 32 0
-- Retrieval info: CONNECT: @data 1 69 32 0 data69x 0 0 32 0
-- Retrieval info: CONNECT: @data 1 6 32 0 data6x 0 0 32 0
-- Retrieval info: CONNECT: @data 1 70 32 0 data70x 0 0 32 0
-- Retrieval info: CONNECT: @data 1 71 32 0 data71x 0 0 32 0
-- Retrieval info: CONNECT: @data 1 72 32 0 data72x 0 0 32 0
-- Retrieval info: CONNECT: @data 1 73 32 0 data73x 0 0 32 0
-- Retrieval info: CONNECT: @data 1 74 32 0 data74x 0 0 32 0
-- Retrieval info: CONNECT: @data 1 75 32 0 data75x 0 0 32 0
-- Retrieval info: CONNECT: @data 1 76 32 0 data76x 0 0 32 0
-- Retrieval info: CONNECT: @data 1 77 32 0 data77x 0 0 32 0
-- Retrieval info: CONNECT: @data 1 78 32 0 data78x 0 0 32 0
-- Retrieval info: CONNECT: @data 1 79 32 0 data79x 0 0 32 0
-- Retrieval info: CONNECT: @data 1 7 32 0 data7x 0 0 32 0
-- Retrieval info: CONNECT: @data 1 80 32 0 data80x 0 0 32 0
-- Retrieval info: CONNECT: @data 1 81 32 0 data81x 0 0 32 0
-- Retrieval info: CONNECT: @data 1 82 32 0 data82x 0 0 32 0
-- Retrieval info: CONNECT: @data 1 83 32 0 data83x 0 0 32 0
-- Retrieval info: CONNECT: @data 1 84 32 0 data84x 0 0 32 0
-- Retrieval info: CONNECT: @data 1 85 32 0 data85x 0 0 32 0
-- Retrieval info: CONNECT: @data 1 86 32 0 data86x 0 0 32 0
-- Retrieval info: CONNECT: @data 1 87 32 0 data87x 0 0 32 0
-- Retrieval info: CONNECT: @data 1 88 32 0 data88x 0 0 32 0
-- Retrieval info: CONNECT: @data 1 89 32 0 data89x 0 0 32 0
-- Retrieval info: CONNECT: @data 1 8 32 0 data8x 0 0 32 0
-- Retrieval info: CONNECT: @data 1 90 32 0 data90x 0 0 32 0
-- Retrieval info: CONNECT: @data 1 91 32 0 data91x 0 0 32 0
-- Retrieval info: CONNECT: @data 1 92 32 0 data92x 0 0 32 0
-- Retrieval info: CONNECT: @data 1 93 32 0 data93x 0 0 32 0
-- Retrieval info: CONNECT: @data 1 94 32 0 data94x 0 0 32 0
-- Retrieval info: CONNECT: @data 1 95 32 0 data95x 0 0 32 0
-- Retrieval info: CONNECT: @data 1 96 32 0 data96x 0 0 32 0
-- Retrieval info: CONNECT: @data 1 97 32 0 data97x 0 0 32 0
-- Retrieval info: CONNECT: @data 1 98 32 0 data98x 0 0 32 0
-- Retrieval info: CONNECT: @data 1 99 32 0 data99x 0 0 32 0
-- Retrieval info: CONNECT: @data 1 9 32 0 data9x 0 0 32 0
-- Retrieval info: CONNECT: @sel 0 0 7 0 sel 0 0 7 0
-- Retrieval info: CONNECT: result 0 0 32 0 @result 0 0 32 0
-- Retrieval info: GEN_FILE: TYPE_NORMAL out_mux.vhd TRUE
-- Retrieval info: GEN_FILE: TYPE_NORMAL out_mux.inc FALSE
-- Retrieval info: GEN_FILE: TYPE_NORMAL out_mux.cmp TRUE
-- Retrieval info: GEN_FILE: TYPE_NORMAL out_mux.bsf FALSE
-- Retrieval info: GEN_FILE: TYPE_NORMAL out_mux_inst.vhd FALSE
-- Retrieval info: LIB_FILE: lpm
