library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity Mux19 is
port(
	U1out,fxs1out: out std_logic_vector(15 downto 0);
	regin: in std_logic_vector(15 downto 0);
	ctrl: in std_logic_vector(1 downto 0)
	);
end Mux19;

architecture bhv of Mux19 is
begin
	process(ctrl,regin)

	variable outTemp : std_logic_vector(15 downto 0);
	begin
		if ctrl = "01" then
			U1out <= regin;
		elsif ctrl = "10" then
			fxs1out <= regin;
		
		end if;
		
	end process;
end bhv;