-- megafunction wizard: %LPM_MUX%
-- GENERATION: STANDARD
-- VERSION: WM1.0
-- MODULE: LPM_MUX 

-- ============================================================
-- File Name: AU_MUX.vhd
-- Megafunction Name(s):
-- 			LPM_MUX
--
-- Simulation Library Files(s):
-- 			lpm
-- ============================================================
-- ************************************************************
-- THIS IS A WIZARD-GENERATED FILE. DO NOT EDIT THIS FILE!
--
-- 18.1.0 Build 625 09/12/2018 SJ Lite Edition
-- ************************************************************


--Copyright (C) 2018  Intel Corporation. All rights reserved.
--Your use of Intel Corporation's design tools, logic functions 
--and other software and tools, and its AMPP partner logic 
--functions, and any output files from any of the foregoing 
--(including device programming or simulation files), and any 
--associated documentation or information are expressly subject 
--to the terms and conditions of the Intel Program License 
--Subscription Agreement, the Intel Quartus Prime License Agreement,
--the Intel FPGA IP License Agreement, or other applicable license
--agreement, including, without limitation, that your use is for
--the sole purpose of programming logic devices manufactured by
--Intel and sold by Intel or its authorized distributors.  Please
--refer to the applicable agreement for further details.


LIBRARY ieee;
USE ieee.std_logic_1164.all;

LIBRARY lpm;
USE lpm.lpm_components.all;

ENTITY AU_MUX IS
	PORT
	(
		data0x		: IN STD_LOGIC_VECTOR (1 DOWNTO 0);
		data10x		: IN STD_LOGIC_VECTOR (1 DOWNTO 0);
		data11x		: IN STD_LOGIC_VECTOR (1 DOWNTO 0);
		data12x		: IN STD_LOGIC_VECTOR (1 DOWNTO 0);
		data13x		: IN STD_LOGIC_VECTOR (1 DOWNTO 0);
		data14x		: IN STD_LOGIC_VECTOR (1 DOWNTO 0);
		data15x		: IN STD_LOGIC_VECTOR (1 DOWNTO 0);
		data16x		: IN STD_LOGIC_VECTOR (1 DOWNTO 0);
		data17x		: IN STD_LOGIC_VECTOR (1 DOWNTO 0);
		data18x		: IN STD_LOGIC_VECTOR (1 DOWNTO 0);
		data19x		: IN STD_LOGIC_VECTOR (1 DOWNTO 0);
		data1x		: IN STD_LOGIC_VECTOR (1 DOWNTO 0);
		data20x		: IN STD_LOGIC_VECTOR (1 DOWNTO 0);
		data21x		: IN STD_LOGIC_VECTOR (1 DOWNTO 0);
		data22x		: IN STD_LOGIC_VECTOR (1 DOWNTO 0);
		data23x		: IN STD_LOGIC_VECTOR (1 DOWNTO 0);
		data24x		: IN STD_LOGIC_VECTOR (1 DOWNTO 0);
		data25x		: IN STD_LOGIC_VECTOR (1 DOWNTO 0);
		data26x		: IN STD_LOGIC_VECTOR (1 DOWNTO 0);
		data27x		: IN STD_LOGIC_VECTOR (1 DOWNTO 0);
		data28x		: IN STD_LOGIC_VECTOR (1 DOWNTO 0);
		data29x		: IN STD_LOGIC_VECTOR (1 DOWNTO 0);
		data2x		: IN STD_LOGIC_VECTOR (1 DOWNTO 0);
		data30x		: IN STD_LOGIC_VECTOR (1 DOWNTO 0);
		data31x		: IN STD_LOGIC_VECTOR (1 DOWNTO 0);
		data32x		: IN STD_LOGIC_VECTOR (1 DOWNTO 0);
		data33x		: IN STD_LOGIC_VECTOR (1 DOWNTO 0);
		data34x		: IN STD_LOGIC_VECTOR (1 DOWNTO 0);
		data35x		: IN STD_LOGIC_VECTOR (1 DOWNTO 0);
		data36x		: IN STD_LOGIC_VECTOR (1 DOWNTO 0);
		data37x		: IN STD_LOGIC_VECTOR (1 DOWNTO 0);
		data38x		: IN STD_LOGIC_VECTOR (1 DOWNTO 0);
		data39x		: IN STD_LOGIC_VECTOR (1 DOWNTO 0);
		data3x		: IN STD_LOGIC_VECTOR (1 DOWNTO 0);
		data40x		: IN STD_LOGIC_VECTOR (1 DOWNTO 0);
		data41x		: IN STD_LOGIC_VECTOR (1 DOWNTO 0);
		data42x		: IN STD_LOGIC_VECTOR (1 DOWNTO 0);
		data43x		: IN STD_LOGIC_VECTOR (1 DOWNTO 0);
		data44x		: IN STD_LOGIC_VECTOR (1 DOWNTO 0);
		data45x		: IN STD_LOGIC_VECTOR (1 DOWNTO 0);
		data46x		: IN STD_LOGIC_VECTOR (1 DOWNTO 0);
		data47x		: IN STD_LOGIC_VECTOR (1 DOWNTO 0);
		data48x		: IN STD_LOGIC_VECTOR (1 DOWNTO 0);
		data49x		: IN STD_LOGIC_VECTOR (1 DOWNTO 0);
		data4x		: IN STD_LOGIC_VECTOR (1 DOWNTO 0);
		data50x		: IN STD_LOGIC_VECTOR (1 DOWNTO 0);
		data51x		: IN STD_LOGIC_VECTOR (1 DOWNTO 0);
		data52x		: IN STD_LOGIC_VECTOR (1 DOWNTO 0);
		data53x		: IN STD_LOGIC_VECTOR (1 DOWNTO 0);
		data54x		: IN STD_LOGIC_VECTOR (1 DOWNTO 0);
		data55x		: IN STD_LOGIC_VECTOR (1 DOWNTO 0);
		data56x		: IN STD_LOGIC_VECTOR (1 DOWNTO 0);
		data57x		: IN STD_LOGIC_VECTOR (1 DOWNTO 0);
		data58x		: IN STD_LOGIC_VECTOR (1 DOWNTO 0);
		data59x		: IN STD_LOGIC_VECTOR (1 DOWNTO 0);
		data5x		: IN STD_LOGIC_VECTOR (1 DOWNTO 0);
		data60x		: IN STD_LOGIC_VECTOR (1 DOWNTO 0);
		data61x		: IN STD_LOGIC_VECTOR (1 DOWNTO 0);
		data62x		: IN STD_LOGIC_VECTOR (1 DOWNTO 0);
		data63x		: IN STD_LOGIC_VECTOR (1 DOWNTO 0);
		data6x		: IN STD_LOGIC_VECTOR (1 DOWNTO 0);
		data7x		: IN STD_LOGIC_VECTOR (1 DOWNTO 0);
		data8x		: IN STD_LOGIC_VECTOR (1 DOWNTO 0);
		data9x		: IN STD_LOGIC_VECTOR (1 DOWNTO 0);
		sel		: IN STD_LOGIC_VECTOR (5 DOWNTO 0);
		result		: OUT STD_LOGIC_VECTOR (1 DOWNTO 0)
	);
END AU_MUX;


ARCHITECTURE SYN OF au_mux IS

--	type STD_LOGIC_2D is array (NATURAL RANGE <>, NATURAL RANGE <>) of STD_LOGIC;

	SIGNAL sub_wire0	: STD_LOGIC_VECTOR (1 DOWNTO 0);
	SIGNAL sub_wire1	: STD_LOGIC_2D (63 DOWNTO 0, 1 DOWNTO 0);
	SIGNAL sub_wire2	: STD_LOGIC_VECTOR (1 DOWNTO 0);
	SIGNAL sub_wire3	: STD_LOGIC_VECTOR (1 DOWNTO 0);
	SIGNAL sub_wire4	: STD_LOGIC_VECTOR (1 DOWNTO 0);
	SIGNAL sub_wire5	: STD_LOGIC_VECTOR (1 DOWNTO 0);
	SIGNAL sub_wire6	: STD_LOGIC_VECTOR (1 DOWNTO 0);
	SIGNAL sub_wire7	: STD_LOGIC_VECTOR (1 DOWNTO 0);
	SIGNAL sub_wire8	: STD_LOGIC_VECTOR (1 DOWNTO 0);
	SIGNAL sub_wire9	: STD_LOGIC_VECTOR (1 DOWNTO 0);
	SIGNAL sub_wire10	: STD_LOGIC_VECTOR (1 DOWNTO 0);
	SIGNAL sub_wire11	: STD_LOGIC_VECTOR (1 DOWNTO 0);
	SIGNAL sub_wire12	: STD_LOGIC_VECTOR (1 DOWNTO 0);
	SIGNAL sub_wire13	: STD_LOGIC_VECTOR (1 DOWNTO 0);
	SIGNAL sub_wire14	: STD_LOGIC_VECTOR (1 DOWNTO 0);
	SIGNAL sub_wire15	: STD_LOGIC_VECTOR (1 DOWNTO 0);
	SIGNAL sub_wire16	: STD_LOGIC_VECTOR (1 DOWNTO 0);
	SIGNAL sub_wire17	: STD_LOGIC_VECTOR (1 DOWNTO 0);
	SIGNAL sub_wire18	: STD_LOGIC_VECTOR (1 DOWNTO 0);
	SIGNAL sub_wire19	: STD_LOGIC_VECTOR (1 DOWNTO 0);
	SIGNAL sub_wire20	: STD_LOGIC_VECTOR (1 DOWNTO 0);
	SIGNAL sub_wire21	: STD_LOGIC_VECTOR (1 DOWNTO 0);
	SIGNAL sub_wire22	: STD_LOGIC_VECTOR (1 DOWNTO 0);
	SIGNAL sub_wire23	: STD_LOGIC_VECTOR (1 DOWNTO 0);
	SIGNAL sub_wire24	: STD_LOGIC_VECTOR (1 DOWNTO 0);
	SIGNAL sub_wire25	: STD_LOGIC_VECTOR (1 DOWNTO 0);
	SIGNAL sub_wire26	: STD_LOGIC_VECTOR (1 DOWNTO 0);
	SIGNAL sub_wire27	: STD_LOGIC_VECTOR (1 DOWNTO 0);
	SIGNAL sub_wire28	: STD_LOGIC_VECTOR (1 DOWNTO 0);
	SIGNAL sub_wire29	: STD_LOGIC_VECTOR (1 DOWNTO 0);
	SIGNAL sub_wire30	: STD_LOGIC_VECTOR (1 DOWNTO 0);
	SIGNAL sub_wire31	: STD_LOGIC_VECTOR (1 DOWNTO 0);
	SIGNAL sub_wire32	: STD_LOGIC_VECTOR (1 DOWNTO 0);
	SIGNAL sub_wire33	: STD_LOGIC_VECTOR (1 DOWNTO 0);
	SIGNAL sub_wire34	: STD_LOGIC_VECTOR (1 DOWNTO 0);
	SIGNAL sub_wire35	: STD_LOGIC_VECTOR (1 DOWNTO 0);
	SIGNAL sub_wire36	: STD_LOGIC_VECTOR (1 DOWNTO 0);
	SIGNAL sub_wire37	: STD_LOGIC_VECTOR (1 DOWNTO 0);
	SIGNAL sub_wire38	: STD_LOGIC_VECTOR (1 DOWNTO 0);
	SIGNAL sub_wire39	: STD_LOGIC_VECTOR (1 DOWNTO 0);
	SIGNAL sub_wire40	: STD_LOGIC_VECTOR (1 DOWNTO 0);
	SIGNAL sub_wire41	: STD_LOGIC_VECTOR (1 DOWNTO 0);
	SIGNAL sub_wire42	: STD_LOGIC_VECTOR (1 DOWNTO 0);
	SIGNAL sub_wire43	: STD_LOGIC_VECTOR (1 DOWNTO 0);
	SIGNAL sub_wire44	: STD_LOGIC_VECTOR (1 DOWNTO 0);
	SIGNAL sub_wire45	: STD_LOGIC_VECTOR (1 DOWNTO 0);
	SIGNAL sub_wire46	: STD_LOGIC_VECTOR (1 DOWNTO 0);
	SIGNAL sub_wire47	: STD_LOGIC_VECTOR (1 DOWNTO 0);
	SIGNAL sub_wire48	: STD_LOGIC_VECTOR (1 DOWNTO 0);
	SIGNAL sub_wire49	: STD_LOGIC_VECTOR (1 DOWNTO 0);
	SIGNAL sub_wire50	: STD_LOGIC_VECTOR (1 DOWNTO 0);
	SIGNAL sub_wire51	: STD_LOGIC_VECTOR (1 DOWNTO 0);
	SIGNAL sub_wire52	: STD_LOGIC_VECTOR (1 DOWNTO 0);
	SIGNAL sub_wire53	: STD_LOGIC_VECTOR (1 DOWNTO 0);
	SIGNAL sub_wire54	: STD_LOGIC_VECTOR (1 DOWNTO 0);
	SIGNAL sub_wire55	: STD_LOGIC_VECTOR (1 DOWNTO 0);
	SIGNAL sub_wire56	: STD_LOGIC_VECTOR (1 DOWNTO 0);
	SIGNAL sub_wire57	: STD_LOGIC_VECTOR (1 DOWNTO 0);
	SIGNAL sub_wire58	: STD_LOGIC_VECTOR (1 DOWNTO 0);
	SIGNAL sub_wire59	: STD_LOGIC_VECTOR (1 DOWNTO 0);
	SIGNAL sub_wire60	: STD_LOGIC_VECTOR (1 DOWNTO 0);
	SIGNAL sub_wire61	: STD_LOGIC_VECTOR (1 DOWNTO 0);
	SIGNAL sub_wire62	: STD_LOGIC_VECTOR (1 DOWNTO 0);
	SIGNAL sub_wire63	: STD_LOGIC_VECTOR (1 DOWNTO 0);
	SIGNAL sub_wire64	: STD_LOGIC_VECTOR (1 DOWNTO 0);
	SIGNAL sub_wire65	: STD_LOGIC_VECTOR (1 DOWNTO 0);

BEGIN
	sub_wire64    <= data0x(1 DOWNTO 0);
	sub_wire63    <= data1x(1 DOWNTO 0);
	sub_wire62    <= data2x(1 DOWNTO 0);
	sub_wire61    <= data3x(1 DOWNTO 0);
	sub_wire60    <= data4x(1 DOWNTO 0);
	sub_wire59    <= data5x(1 DOWNTO 0);
	sub_wire58    <= data6x(1 DOWNTO 0);
	sub_wire57    <= data7x(1 DOWNTO 0);
	sub_wire56    <= data8x(1 DOWNTO 0);
	sub_wire55    <= data9x(1 DOWNTO 0);
	sub_wire54    <= data10x(1 DOWNTO 0);
	sub_wire53    <= data11x(1 DOWNTO 0);
	sub_wire52    <= data12x(1 DOWNTO 0);
	sub_wire51    <= data13x(1 DOWNTO 0);
	sub_wire50    <= data14x(1 DOWNTO 0);
	sub_wire49    <= data15x(1 DOWNTO 0);
	sub_wire48    <= data16x(1 DOWNTO 0);
	sub_wire47    <= data17x(1 DOWNTO 0);
	sub_wire46    <= data18x(1 DOWNTO 0);
	sub_wire45    <= data19x(1 DOWNTO 0);
	sub_wire44    <= data20x(1 DOWNTO 0);
	sub_wire43    <= data21x(1 DOWNTO 0);
	sub_wire42    <= data22x(1 DOWNTO 0);
	sub_wire41    <= data23x(1 DOWNTO 0);
	sub_wire40    <= data24x(1 DOWNTO 0);
	sub_wire39    <= data25x(1 DOWNTO 0);
	sub_wire38    <= data26x(1 DOWNTO 0);
	sub_wire37    <= data27x(1 DOWNTO 0);
	sub_wire36    <= data28x(1 DOWNTO 0);
	sub_wire35    <= data29x(1 DOWNTO 0);
	sub_wire34    <= data30x(1 DOWNTO 0);
	sub_wire33    <= data31x(1 DOWNTO 0);
	sub_wire32    <= data32x(1 DOWNTO 0);
	sub_wire31    <= data33x(1 DOWNTO 0);
	sub_wire30    <= data34x(1 DOWNTO 0);
	sub_wire29    <= data35x(1 DOWNTO 0);
	sub_wire28    <= data36x(1 DOWNTO 0);
	sub_wire27    <= data37x(1 DOWNTO 0);
	sub_wire26    <= data38x(1 DOWNTO 0);
	sub_wire25    <= data39x(1 DOWNTO 0);
	sub_wire24    <= data40x(1 DOWNTO 0);
	sub_wire23    <= data41x(1 DOWNTO 0);
	sub_wire22    <= data42x(1 DOWNTO 0);
	sub_wire21    <= data43x(1 DOWNTO 0);
	sub_wire20    <= data44x(1 DOWNTO 0);
	sub_wire19    <= data45x(1 DOWNTO 0);
	sub_wire18    <= data46x(1 DOWNTO 0);
	sub_wire17    <= data47x(1 DOWNTO 0);
	sub_wire16    <= data48x(1 DOWNTO 0);
	sub_wire15    <= data49x(1 DOWNTO 0);
	sub_wire14    <= data50x(1 DOWNTO 0);
	sub_wire13    <= data51x(1 DOWNTO 0);
	sub_wire12    <= data52x(1 DOWNTO 0);
	sub_wire11    <= data53x(1 DOWNTO 0);
	sub_wire10    <= data54x(1 DOWNTO 0);
	sub_wire9    <= data55x(1 DOWNTO 0);
	sub_wire8    <= data56x(1 DOWNTO 0);
	sub_wire7    <= data57x(1 DOWNTO 0);
	sub_wire6    <= data58x(1 DOWNTO 0);
	sub_wire5    <= data59x(1 DOWNTO 0);
	sub_wire4    <= data60x(1 DOWNTO 0);
	sub_wire3    <= data61x(1 DOWNTO 0);
	sub_wire2    <= data62x(1 DOWNTO 0);
	sub_wire0    <= data63x(1 DOWNTO 0);
	sub_wire1(63, 0)    <= sub_wire0(0);
	sub_wire1(63, 1)    <= sub_wire0(1);
	sub_wire1(62, 0)    <= sub_wire2(0);
	sub_wire1(62, 1)    <= sub_wire2(1);
	sub_wire1(61, 0)    <= sub_wire3(0);
	sub_wire1(61, 1)    <= sub_wire3(1);
	sub_wire1(60, 0)    <= sub_wire4(0);
	sub_wire1(60, 1)    <= sub_wire4(1);
	sub_wire1(59, 0)    <= sub_wire5(0);
	sub_wire1(59, 1)    <= sub_wire5(1);
	sub_wire1(58, 0)    <= sub_wire6(0);
	sub_wire1(58, 1)    <= sub_wire6(1);
	sub_wire1(57, 0)    <= sub_wire7(0);
	sub_wire1(57, 1)    <= sub_wire7(1);
	sub_wire1(56, 0)    <= sub_wire8(0);
	sub_wire1(56, 1)    <= sub_wire8(1);
	sub_wire1(55, 0)    <= sub_wire9(0);
	sub_wire1(55, 1)    <= sub_wire9(1);
	sub_wire1(54, 0)    <= sub_wire10(0);
	sub_wire1(54, 1)    <= sub_wire10(1);
	sub_wire1(53, 0)    <= sub_wire11(0);
	sub_wire1(53, 1)    <= sub_wire11(1);
	sub_wire1(52, 0)    <= sub_wire12(0);
	sub_wire1(52, 1)    <= sub_wire12(1);
	sub_wire1(51, 0)    <= sub_wire13(0);
	sub_wire1(51, 1)    <= sub_wire13(1);
	sub_wire1(50, 0)    <= sub_wire14(0);
	sub_wire1(50, 1)    <= sub_wire14(1);
	sub_wire1(49, 0)    <= sub_wire15(0);
	sub_wire1(49, 1)    <= sub_wire15(1);
	sub_wire1(48, 0)    <= sub_wire16(0);
	sub_wire1(48, 1)    <= sub_wire16(1);
	sub_wire1(47, 0)    <= sub_wire17(0);
	sub_wire1(47, 1)    <= sub_wire17(1);
	sub_wire1(46, 0)    <= sub_wire18(0);
	sub_wire1(46, 1)    <= sub_wire18(1);
	sub_wire1(45, 0)    <= sub_wire19(0);
	sub_wire1(45, 1)    <= sub_wire19(1);
	sub_wire1(44, 0)    <= sub_wire20(0);
	sub_wire1(44, 1)    <= sub_wire20(1);
	sub_wire1(43, 0)    <= sub_wire21(0);
	sub_wire1(43, 1)    <= sub_wire21(1);
	sub_wire1(42, 0)    <= sub_wire22(0);
	sub_wire1(42, 1)    <= sub_wire22(1);
	sub_wire1(41, 0)    <= sub_wire23(0);
	sub_wire1(41, 1)    <= sub_wire23(1);
	sub_wire1(40, 0)    <= sub_wire24(0);
	sub_wire1(40, 1)    <= sub_wire24(1);
	sub_wire1(39, 0)    <= sub_wire25(0);
	sub_wire1(39, 1)    <= sub_wire25(1);
	sub_wire1(38, 0)    <= sub_wire26(0);
	sub_wire1(38, 1)    <= sub_wire26(1);
	sub_wire1(37, 0)    <= sub_wire27(0);
	sub_wire1(37, 1)    <= sub_wire27(1);
	sub_wire1(36, 0)    <= sub_wire28(0);
	sub_wire1(36, 1)    <= sub_wire28(1);
	sub_wire1(35, 0)    <= sub_wire29(0);
	sub_wire1(35, 1)    <= sub_wire29(1);
	sub_wire1(34, 0)    <= sub_wire30(0);
	sub_wire1(34, 1)    <= sub_wire30(1);
	sub_wire1(33, 0)    <= sub_wire31(0);
	sub_wire1(33, 1)    <= sub_wire31(1);
	sub_wire1(32, 0)    <= sub_wire32(0);
	sub_wire1(32, 1)    <= sub_wire32(1);
	sub_wire1(31, 0)    <= sub_wire33(0);
	sub_wire1(31, 1)    <= sub_wire33(1);
	sub_wire1(30, 0)    <= sub_wire34(0);
	sub_wire1(30, 1)    <= sub_wire34(1);
	sub_wire1(29, 0)    <= sub_wire35(0);
	sub_wire1(29, 1)    <= sub_wire35(1);
	sub_wire1(28, 0)    <= sub_wire36(0);
	sub_wire1(28, 1)    <= sub_wire36(1);
	sub_wire1(27, 0)    <= sub_wire37(0);
	sub_wire1(27, 1)    <= sub_wire37(1);
	sub_wire1(26, 0)    <= sub_wire38(0);
	sub_wire1(26, 1)    <= sub_wire38(1);
	sub_wire1(25, 0)    <= sub_wire39(0);
	sub_wire1(25, 1)    <= sub_wire39(1);
	sub_wire1(24, 0)    <= sub_wire40(0);
	sub_wire1(24, 1)    <= sub_wire40(1);
	sub_wire1(23, 0)    <= sub_wire41(0);
	sub_wire1(23, 1)    <= sub_wire41(1);
	sub_wire1(22, 0)    <= sub_wire42(0);
	sub_wire1(22, 1)    <= sub_wire42(1);
	sub_wire1(21, 0)    <= sub_wire43(0);
	sub_wire1(21, 1)    <= sub_wire43(1);
	sub_wire1(20, 0)    <= sub_wire44(0);
	sub_wire1(20, 1)    <= sub_wire44(1);
	sub_wire1(19, 0)    <= sub_wire45(0);
	sub_wire1(19, 1)    <= sub_wire45(1);
	sub_wire1(18, 0)    <= sub_wire46(0);
	sub_wire1(18, 1)    <= sub_wire46(1);
	sub_wire1(17, 0)    <= sub_wire47(0);
	sub_wire1(17, 1)    <= sub_wire47(1);
	sub_wire1(16, 0)    <= sub_wire48(0);
	sub_wire1(16, 1)    <= sub_wire48(1);
	sub_wire1(15, 0)    <= sub_wire49(0);
	sub_wire1(15, 1)    <= sub_wire49(1);
	sub_wire1(14, 0)    <= sub_wire50(0);
	sub_wire1(14, 1)    <= sub_wire50(1);
	sub_wire1(13, 0)    <= sub_wire51(0);
	sub_wire1(13, 1)    <= sub_wire51(1);
	sub_wire1(12, 0)    <= sub_wire52(0);
	sub_wire1(12, 1)    <= sub_wire52(1);
	sub_wire1(11, 0)    <= sub_wire53(0);
	sub_wire1(11, 1)    <= sub_wire53(1);
	sub_wire1(10, 0)    <= sub_wire54(0);
	sub_wire1(10, 1)    <= sub_wire54(1);
	sub_wire1(9, 0)    <= sub_wire55(0);
	sub_wire1(9, 1)    <= sub_wire55(1);
	sub_wire1(8, 0)    <= sub_wire56(0);
	sub_wire1(8, 1)    <= sub_wire56(1);
	sub_wire1(7, 0)    <= sub_wire57(0);
	sub_wire1(7, 1)    <= sub_wire57(1);
	sub_wire1(6, 0)    <= sub_wire58(0);
	sub_wire1(6, 1)    <= sub_wire58(1);
	sub_wire1(5, 0)    <= sub_wire59(0);
	sub_wire1(5, 1)    <= sub_wire59(1);
	sub_wire1(4, 0)    <= sub_wire60(0);
	sub_wire1(4, 1)    <= sub_wire60(1);
	sub_wire1(3, 0)    <= sub_wire61(0);
	sub_wire1(3, 1)    <= sub_wire61(1);
	sub_wire1(2, 0)    <= sub_wire62(0);
	sub_wire1(2, 1)    <= sub_wire62(1);
	sub_wire1(1, 0)    <= sub_wire63(0);
	sub_wire1(1, 1)    <= sub_wire63(1);
	sub_wire1(0, 0)    <= sub_wire64(0);
	sub_wire1(0, 1)    <= sub_wire64(1);
	result    <= sub_wire65(1 DOWNTO 0);

	LPM_MUX_component : LPM_MUX
	GENERIC MAP (
		lpm_size => 64,
		lpm_type => "LPM_MUX",
		lpm_width => 2,
		lpm_widths => 6
	)
	PORT MAP (
		data => sub_wire1,
		sel => sel,
		result => sub_wire65
	);



END SYN;

-- ============================================================
-- CNX file retrieval info
-- ============================================================
-- Retrieval info: PRIVATE: INTENDED_DEVICE_FAMILY STRING "Cyclone IV E"
-- Retrieval info: PRIVATE: SYNTH_WRAPPER_GEN_POSTFIX STRING "0"
-- Retrieval info: PRIVATE: new_diagram STRING "1"
-- Retrieval info: LIBRARY: lpm lpm.lpm_components.all
-- Retrieval info: CONSTANT: LPM_SIZE NUMERIC "64"
-- Retrieval info: CONSTANT: LPM_TYPE STRING "LPM_MUX"
-- Retrieval info: CONSTANT: LPM_WIDTH NUMERIC "2"
-- Retrieval info: CONSTANT: LPM_WIDTHS NUMERIC "6"
-- Retrieval info: USED_PORT: data0x 0 0 2 0 INPUT NODEFVAL "data0x[1..0]"
-- Retrieval info: USED_PORT: data10x 0 0 2 0 INPUT NODEFVAL "data10x[1..0]"
-- Retrieval info: USED_PORT: data11x 0 0 2 0 INPUT NODEFVAL "data11x[1..0]"
-- Retrieval info: USED_PORT: data12x 0 0 2 0 INPUT NODEFVAL "data12x[1..0]"
-- Retrieval info: USED_PORT: data13x 0 0 2 0 INPUT NODEFVAL "data13x[1..0]"
-- Retrieval info: USED_PORT: data14x 0 0 2 0 INPUT NODEFVAL "data14x[1..0]"
-- Retrieval info: USED_PORT: data15x 0 0 2 0 INPUT NODEFVAL "data15x[1..0]"
-- Retrieval info: USED_PORT: data16x 0 0 2 0 INPUT NODEFVAL "data16x[1..0]"
-- Retrieval info: USED_PORT: data17x 0 0 2 0 INPUT NODEFVAL "data17x[1..0]"
-- Retrieval info: USED_PORT: data18x 0 0 2 0 INPUT NODEFVAL "data18x[1..0]"
-- Retrieval info: USED_PORT: data19x 0 0 2 0 INPUT NODEFVAL "data19x[1..0]"
-- Retrieval info: USED_PORT: data1x 0 0 2 0 INPUT NODEFVAL "data1x[1..0]"
-- Retrieval info: USED_PORT: data20x 0 0 2 0 INPUT NODEFVAL "data20x[1..0]"
-- Retrieval info: USED_PORT: data21x 0 0 2 0 INPUT NODEFVAL "data21x[1..0]"
-- Retrieval info: USED_PORT: data22x 0 0 2 0 INPUT NODEFVAL "data22x[1..0]"
-- Retrieval info: USED_PORT: data23x 0 0 2 0 INPUT NODEFVAL "data23x[1..0]"
-- Retrieval info: USED_PORT: data24x 0 0 2 0 INPUT NODEFVAL "data24x[1..0]"
-- Retrieval info: USED_PORT: data25x 0 0 2 0 INPUT NODEFVAL "data25x[1..0]"
-- Retrieval info: USED_PORT: data26x 0 0 2 0 INPUT NODEFVAL "data26x[1..0]"
-- Retrieval info: USED_PORT: data27x 0 0 2 0 INPUT NODEFVAL "data27x[1..0]"
-- Retrieval info: USED_PORT: data28x 0 0 2 0 INPUT NODEFVAL "data28x[1..0]"
-- Retrieval info: USED_PORT: data29x 0 0 2 0 INPUT NODEFVAL "data29x[1..0]"
-- Retrieval info: USED_PORT: data2x 0 0 2 0 INPUT NODEFVAL "data2x[1..0]"
-- Retrieval info: USED_PORT: data30x 0 0 2 0 INPUT NODEFVAL "data30x[1..0]"
-- Retrieval info: USED_PORT: data31x 0 0 2 0 INPUT NODEFVAL "data31x[1..0]"
-- Retrieval info: USED_PORT: data32x 0 0 2 0 INPUT NODEFVAL "data32x[1..0]"
-- Retrieval info: USED_PORT: data33x 0 0 2 0 INPUT NODEFVAL "data33x[1..0]"
-- Retrieval info: USED_PORT: data34x 0 0 2 0 INPUT NODEFVAL "data34x[1..0]"
-- Retrieval info: USED_PORT: data35x 0 0 2 0 INPUT NODEFVAL "data35x[1..0]"
-- Retrieval info: USED_PORT: data36x 0 0 2 0 INPUT NODEFVAL "data36x[1..0]"
-- Retrieval info: USED_PORT: data37x 0 0 2 0 INPUT NODEFVAL "data37x[1..0]"
-- Retrieval info: USED_PORT: data38x 0 0 2 0 INPUT NODEFVAL "data38x[1..0]"
-- Retrieval info: USED_PORT: data39x 0 0 2 0 INPUT NODEFVAL "data39x[1..0]"
-- Retrieval info: USED_PORT: data3x 0 0 2 0 INPUT NODEFVAL "data3x[1..0]"
-- Retrieval info: USED_PORT: data40x 0 0 2 0 INPUT NODEFVAL "data40x[1..0]"
-- Retrieval info: USED_PORT: data41x 0 0 2 0 INPUT NODEFVAL "data41x[1..0]"
-- Retrieval info: USED_PORT: data42x 0 0 2 0 INPUT NODEFVAL "data42x[1..0]"
-- Retrieval info: USED_PORT: data43x 0 0 2 0 INPUT NODEFVAL "data43x[1..0]"
-- Retrieval info: USED_PORT: data44x 0 0 2 0 INPUT NODEFVAL "data44x[1..0]"
-- Retrieval info: USED_PORT: data45x 0 0 2 0 INPUT NODEFVAL "data45x[1..0]"
-- Retrieval info: USED_PORT: data46x 0 0 2 0 INPUT NODEFVAL "data46x[1..0]"
-- Retrieval info: USED_PORT: data47x 0 0 2 0 INPUT NODEFVAL "data47x[1..0]"
-- Retrieval info: USED_PORT: data48x 0 0 2 0 INPUT NODEFVAL "data48x[1..0]"
-- Retrieval info: USED_PORT: data49x 0 0 2 0 INPUT NODEFVAL "data49x[1..0]"
-- Retrieval info: USED_PORT: data4x 0 0 2 0 INPUT NODEFVAL "data4x[1..0]"
-- Retrieval info: USED_PORT: data50x 0 0 2 0 INPUT NODEFVAL "data50x[1..0]"
-- Retrieval info: USED_PORT: data51x 0 0 2 0 INPUT NODEFVAL "data51x[1..0]"
-- Retrieval info: USED_PORT: data52x 0 0 2 0 INPUT NODEFVAL "data52x[1..0]"
-- Retrieval info: USED_PORT: data53x 0 0 2 0 INPUT NODEFVAL "data53x[1..0]"
-- Retrieval info: USED_PORT: data54x 0 0 2 0 INPUT NODEFVAL "data54x[1..0]"
-- Retrieval info: USED_PORT: data55x 0 0 2 0 INPUT NODEFVAL "data55x[1..0]"
-- Retrieval info: USED_PORT: data56x 0 0 2 0 INPUT NODEFVAL "data56x[1..0]"
-- Retrieval info: USED_PORT: data57x 0 0 2 0 INPUT NODEFVAL "data57x[1..0]"
-- Retrieval info: USED_PORT: data58x 0 0 2 0 INPUT NODEFVAL "data58x[1..0]"
-- Retrieval info: USED_PORT: data59x 0 0 2 0 INPUT NODEFVAL "data59x[1..0]"
-- Retrieval info: USED_PORT: data5x 0 0 2 0 INPUT NODEFVAL "data5x[1..0]"
-- Retrieval info: USED_PORT: data60x 0 0 2 0 INPUT NODEFVAL "data60x[1..0]"
-- Retrieval info: USED_PORT: data61x 0 0 2 0 INPUT NODEFVAL "data61x[1..0]"
-- Retrieval info: USED_PORT: data62x 0 0 2 0 INPUT NODEFVAL "data62x[1..0]"
-- Retrieval info: USED_PORT: data63x 0 0 2 0 INPUT NODEFVAL "data63x[1..0]"
-- Retrieval info: USED_PORT: data6x 0 0 2 0 INPUT NODEFVAL "data6x[1..0]"
-- Retrieval info: USED_PORT: data7x 0 0 2 0 INPUT NODEFVAL "data7x[1..0]"
-- Retrieval info: USED_PORT: data8x 0 0 2 0 INPUT NODEFVAL "data8x[1..0]"
-- Retrieval info: USED_PORT: data9x 0 0 2 0 INPUT NODEFVAL "data9x[1..0]"
-- Retrieval info: USED_PORT: result 0 0 2 0 OUTPUT NODEFVAL "result[1..0]"
-- Retrieval info: USED_PORT: sel 0 0 6 0 INPUT NODEFVAL "sel[5..0]"
-- Retrieval info: CONNECT: @data 1 0 2 0 data0x 0 0 2 0
-- Retrieval info: CONNECT: @data 1 10 2 0 data10x 0 0 2 0
-- Retrieval info: CONNECT: @data 1 11 2 0 data11x 0 0 2 0
-- Retrieval info: CONNECT: @data 1 12 2 0 data12x 0 0 2 0
-- Retrieval info: CONNECT: @data 1 13 2 0 data13x 0 0 2 0
-- Retrieval info: CONNECT: @data 1 14 2 0 data14x 0 0 2 0
-- Retrieval info: CONNECT: @data 1 15 2 0 data15x 0 0 2 0
-- Retrieval info: CONNECT: @data 1 16 2 0 data16x 0 0 2 0
-- Retrieval info: CONNECT: @data 1 17 2 0 data17x 0 0 2 0
-- Retrieval info: CONNECT: @data 1 18 2 0 data18x 0 0 2 0
-- Retrieval info: CONNECT: @data 1 19 2 0 data19x 0 0 2 0
-- Retrieval info: CONNECT: @data 1 1 2 0 data1x 0 0 2 0
-- Retrieval info: CONNECT: @data 1 20 2 0 data20x 0 0 2 0
-- Retrieval info: CONNECT: @data 1 21 2 0 data21x 0 0 2 0
-- Retrieval info: CONNECT: @data 1 22 2 0 data22x 0 0 2 0
-- Retrieval info: CONNECT: @data 1 23 2 0 data23x 0 0 2 0
-- Retrieval info: CONNECT: @data 1 24 2 0 data24x 0 0 2 0
-- Retrieval info: CONNECT: @data 1 25 2 0 data25x 0 0 2 0
-- Retrieval info: CONNECT: @data 1 26 2 0 data26x 0 0 2 0
-- Retrieval info: CONNECT: @data 1 27 2 0 data27x 0 0 2 0
-- Retrieval info: CONNECT: @data 1 28 2 0 data28x 0 0 2 0
-- Retrieval info: CONNECT: @data 1 29 2 0 data29x 0 0 2 0
-- Retrieval info: CONNECT: @data 1 2 2 0 data2x 0 0 2 0
-- Retrieval info: CONNECT: @data 1 30 2 0 data30x 0 0 2 0
-- Retrieval info: CONNECT: @data 1 31 2 0 data31x 0 0 2 0
-- Retrieval info: CONNECT: @data 1 32 2 0 data32x 0 0 2 0
-- Retrieval info: CONNECT: @data 1 33 2 0 data33x 0 0 2 0
-- Retrieval info: CONNECT: @data 1 34 2 0 data34x 0 0 2 0
-- Retrieval info: CONNECT: @data 1 35 2 0 data35x 0 0 2 0
-- Retrieval info: CONNECT: @data 1 36 2 0 data36x 0 0 2 0
-- Retrieval info: CONNECT: @data 1 37 2 0 data37x 0 0 2 0
-- Retrieval info: CONNECT: @data 1 38 2 0 data38x 0 0 2 0
-- Retrieval info: CONNECT: @data 1 39 2 0 data39x 0 0 2 0
-- Retrieval info: CONNECT: @data 1 3 2 0 data3x 0 0 2 0
-- Retrieval info: CONNECT: @data 1 40 2 0 data40x 0 0 2 0
-- Retrieval info: CONNECT: @data 1 41 2 0 data41x 0 0 2 0
-- Retrieval info: CONNECT: @data 1 42 2 0 data42x 0 0 2 0
-- Retrieval info: CONNECT: @data 1 43 2 0 data43x 0 0 2 0
-- Retrieval info: CONNECT: @data 1 44 2 0 data44x 0 0 2 0
-- Retrieval info: CONNECT: @data 1 45 2 0 data45x 0 0 2 0
-- Retrieval info: CONNECT: @data 1 46 2 0 data46x 0 0 2 0
-- Retrieval info: CONNECT: @data 1 47 2 0 data47x 0 0 2 0
-- Retrieval info: CONNECT: @data 1 48 2 0 data48x 0 0 2 0
-- Retrieval info: CONNECT: @data 1 49 2 0 data49x 0 0 2 0
-- Retrieval info: CONNECT: @data 1 4 2 0 data4x 0 0 2 0
-- Retrieval info: CONNECT: @data 1 50 2 0 data50x 0 0 2 0
-- Retrieval info: CONNECT: @data 1 51 2 0 data51x 0 0 2 0
-- Retrieval info: CONNECT: @data 1 52 2 0 data52x 0 0 2 0
-- Retrieval info: CONNECT: @data 1 53 2 0 data53x 0 0 2 0
-- Retrieval info: CONNECT: @data 1 54 2 0 data54x 0 0 2 0
-- Retrieval info: CONNECT: @data 1 55 2 0 data55x 0 0 2 0
-- Retrieval info: CONNECT: @data 1 56 2 0 data56x 0 0 2 0
-- Retrieval info: CONNECT: @data 1 57 2 0 data57x 0 0 2 0
-- Retrieval info: CONNECT: @data 1 58 2 0 data58x 0 0 2 0
-- Retrieval info: CONNECT: @data 1 59 2 0 data59x 0 0 2 0
-- Retrieval info: CONNECT: @data 1 5 2 0 data5x 0 0 2 0
-- Retrieval info: CONNECT: @data 1 60 2 0 data60x 0 0 2 0
-- Retrieval info: CONNECT: @data 1 61 2 0 data61x 0 0 2 0
-- Retrieval info: CONNECT: @data 1 62 2 0 data62x 0 0 2 0
-- Retrieval info: CONNECT: @data 1 63 2 0 data63x 0 0 2 0
-- Retrieval info: CONNECT: @data 1 6 2 0 data6x 0 0 2 0
-- Retrieval info: CONNECT: @data 1 7 2 0 data7x 0 0 2 0
-- Retrieval info: CONNECT: @data 1 8 2 0 data8x 0 0 2 0
-- Retrieval info: CONNECT: @data 1 9 2 0 data9x 0 0 2 0
-- Retrieval info: CONNECT: @sel 0 0 6 0 sel 0 0 6 0
-- Retrieval info: CONNECT: result 0 0 2 0 @result 0 0 2 0
-- Retrieval info: GEN_FILE: TYPE_NORMAL AU_MUX.vhd TRUE
-- Retrieval info: GEN_FILE: TYPE_NORMAL AU_MUX.inc FALSE
-- Retrieval info: GEN_FILE: TYPE_NORMAL AU_MUX.cmp TRUE
-- Retrieval info: GEN_FILE: TYPE_NORMAL AU_MUX.bsf FALSE
-- Retrieval info: GEN_FILE: TYPE_NORMAL AU_MUX_inst.vhd TRUE
-- Retrieval info: LIB_FILE: lpm
