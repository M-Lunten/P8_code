AU_MUX_inst : AU_MUX PORT MAP (
		data0x	 => data0x_sig,
		data10x	 => data10x_sig,
		data11x	 => data11x_sig,
		data12x	 => data12x_sig,
		data13x	 => data13x_sig,
		data14x	 => data14x_sig,
		data15x	 => data15x_sig,
		data16x	 => data16x_sig,
		data17x	 => data17x_sig,
		data18x	 => data18x_sig,
		data19x	 => data19x_sig,
		data1x	 => data1x_sig,
		data20x	 => data20x_sig,
		data21x	 => data21x_sig,
		data22x	 => data22x_sig,
		data23x	 => data23x_sig,
		data24x	 => data24x_sig,
		data25x	 => data25x_sig,
		data26x	 => data26x_sig,
		data27x	 => data27x_sig,
		data28x	 => data28x_sig,
		data29x	 => data29x_sig,
		data2x	 => data2x_sig,
		data30x	 => data30x_sig,
		data31x	 => data31x_sig,
		data32x	 => data32x_sig,
		data33x	 => data33x_sig,
		data34x	 => data34x_sig,
		data35x	 => data35x_sig,
		data36x	 => data36x_sig,
		data37x	 => data37x_sig,
		data38x	 => data38x_sig,
		data39x	 => data39x_sig,
		data3x	 => data3x_sig,
		data40x	 => data40x_sig,
		data41x	 => data41x_sig,
		data42x	 => data42x_sig,
		data43x	 => data43x_sig,
		data44x	 => data44x_sig,
		data45x	 => data45x_sig,
		data46x	 => data46x_sig,
		data47x	 => data47x_sig,
		data48x	 => data48x_sig,
		data49x	 => data49x_sig,
		data4x	 => data4x_sig,
		data50x	 => data50x_sig,
		data51x	 => data51x_sig,
		data52x	 => data52x_sig,
		data53x	 => data53x_sig,
		data54x	 => data54x_sig,
		data55x	 => data55x_sig,
		data56x	 => data56x_sig,
		data57x	 => data57x_sig,
		data58x	 => data58x_sig,
		data59x	 => data59x_sig,
		data5x	 => data5x_sig,
		data60x	 => data60x_sig,
		data61x	 => data61x_sig,
		data62x	 => data62x_sig,
		data63x	 => data63x_sig,
		data6x	 => data6x_sig,
		data7x	 => data7x_sig,
		data8x	 => data8x_sig,
		data9x	 => data9x_sig,
		sel	 => sel_sig,
		result	 => result_sig
	);
